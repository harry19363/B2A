`timescale 1ns / 1ps

module A2Bn8(
    input clk_i,
    input rst_ni,
    input i_dvld,
    input i_rvld,
    input [11615:0] i_n,
    input [255:0] i_a,
    output [255:0] o_z,
    output o_dvld
	);


endmodule
