//////////////////////////////////////////////////////////////////////////////////
// Company       : TSU
// Engineer      : 
// 
// Create Date   : 2025-03-06
// File Name     : SecAnd_PINI1_n8k32_1.v
// Project Name  : 
// Design Name   : 
// Description   : 
//                
// 
// Dependencies  : 
// 
// Revision      : 
//                 - V1.0 File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// 
// WARNING: THIS FILE IS AUTOGENERATED
// ANY MANUAL CHANGES WILL BE LOST

`timescale 1ns/1ps
module SecAnd_PINI1_n8k32_1(
    input  wire         clk_i,
    input  wire         rst_ni,
    input  wire         i_dvld,
    input  wire         i_rvld,
    input  wire [895:0] i_n,
    input  wire [255:0] i_x,
    input  wire [255:0] i_y,
    output wire [255:0] o_c,
    output wire         o_dvld);

(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire  vldd1;// synopsys keep_signal_name "vldd1" 
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_0;// synopsys keep_signal_name "xd_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_1;// synopsys keep_signal_name "xd_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_2;// synopsys keep_signal_name "xd_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_3;// synopsys keep_signal_name "xd_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_4;// synopsys keep_signal_name "xd_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_5;// synopsys keep_signal_name "xd_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_6;// synopsys keep_signal_name "xd_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xd_7;// synopsys keep_signal_name "xd_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_0;// synopsys keep_signal_name "yd_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_1;// synopsys keep_signal_name "yd_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_2;// synopsys keep_signal_name "yd_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_3;// synopsys keep_signal_name "yd_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_4;// synopsys keep_signal_name "yd_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_5;// synopsys keep_signal_name "yd_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_6;// synopsys keep_signal_name "yd_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yd_7;// synopsys keep_signal_name "yd_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_0;// synopsys keep_signal_name "r_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_1;// synopsys keep_signal_name "r_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_2;// synopsys keep_signal_name "r_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_3;// synopsys keep_signal_name "r_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_4;// synopsys keep_signal_name "r_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_5;// synopsys keep_signal_name "r_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_6;// synopsys keep_signal_name "r_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_7;// synopsys keep_signal_name "r_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_8;// synopsys keep_signal_name "r_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_9;// synopsys keep_signal_name "r_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_10;// synopsys keep_signal_name "r_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_11;// synopsys keep_signal_name "r_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_12;// synopsys keep_signal_name "r_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_13;// synopsys keep_signal_name "r_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_14;// synopsys keep_signal_name "r_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_15;// synopsys keep_signal_name "r_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_16;// synopsys keep_signal_name "r_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_17;// synopsys keep_signal_name "r_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_18;// synopsys keep_signal_name "r_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_19;// synopsys keep_signal_name "r_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_20;// synopsys keep_signal_name "r_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_21;// synopsys keep_signal_name "r_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_22;// synopsys keep_signal_name "r_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_23;// synopsys keep_signal_name "r_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_24;// synopsys keep_signal_name "r_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_25;// synopsys keep_signal_name "r_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_26;// synopsys keep_signal_name "r_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_27;// synopsys keep_signal_name "r_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_28;// synopsys keep_signal_name "r_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_29;// synopsys keep_signal_name "r_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_30;// synopsys keep_signal_name "r_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_31;// synopsys keep_signal_name "r_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_32;// synopsys keep_signal_name "r_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_33;// synopsys keep_signal_name "r_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_34;// synopsys keep_signal_name "r_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_35;// synopsys keep_signal_name "r_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_36;// synopsys keep_signal_name "r_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_37;// synopsys keep_signal_name "r_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_38;// synopsys keep_signal_name "r_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_39;// synopsys keep_signal_name "r_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_40;// synopsys keep_signal_name "r_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_41;// synopsys keep_signal_name "r_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_42;// synopsys keep_signal_name "r_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_43;// synopsys keep_signal_name "r_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_44;// synopsys keep_signal_name "r_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_45;// synopsys keep_signal_name "r_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_46;// synopsys keep_signal_name "r_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_47;// synopsys keep_signal_name "r_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_48;// synopsys keep_signal_name "r_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_49;// synopsys keep_signal_name "r_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_50;// synopsys keep_signal_name "r_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_51;// synopsys keep_signal_name "r_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_52;// synopsys keep_signal_name "r_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_53;// synopsys keep_signal_name "r_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_54;// synopsys keep_signal_name "r_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] r_55;// synopsys keep_signal_name "r_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_0;// synopsys keep_signal_name "yxn_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_1;// synopsys keep_signal_name "yxn_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_2;// synopsys keep_signal_name "yxn_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_3;// synopsys keep_signal_name "yxn_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_4;// synopsys keep_signal_name "yxn_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_5;// synopsys keep_signal_name "yxn_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_6;// synopsys keep_signal_name "yxn_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_7;// synopsys keep_signal_name "yxn_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_8;// synopsys keep_signal_name "yxn_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_9;// synopsys keep_signal_name "yxn_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_10;// synopsys keep_signal_name "yxn_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_11;// synopsys keep_signal_name "yxn_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_12;// synopsys keep_signal_name "yxn_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_13;// synopsys keep_signal_name "yxn_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_14;// synopsys keep_signal_name "yxn_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_15;// synopsys keep_signal_name "yxn_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_16;// synopsys keep_signal_name "yxn_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_17;// synopsys keep_signal_name "yxn_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_18;// synopsys keep_signal_name "yxn_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_19;// synopsys keep_signal_name "yxn_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_20;// synopsys keep_signal_name "yxn_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_21;// synopsys keep_signal_name "yxn_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_22;// synopsys keep_signal_name "yxn_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_23;// synopsys keep_signal_name "yxn_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_24;// synopsys keep_signal_name "yxn_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_25;// synopsys keep_signal_name "yxn_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_26;// synopsys keep_signal_name "yxn_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_27;// synopsys keep_signal_name "yxn_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_28;// synopsys keep_signal_name "yxn_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_29;// synopsys keep_signal_name "yxn_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_30;// synopsys keep_signal_name "yxn_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_31;// synopsys keep_signal_name "yxn_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_32;// synopsys keep_signal_name "yxn_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_33;// synopsys keep_signal_name "yxn_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_34;// synopsys keep_signal_name "yxn_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_35;// synopsys keep_signal_name "yxn_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_36;// synopsys keep_signal_name "yxn_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_37;// synopsys keep_signal_name "yxn_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_38;// synopsys keep_signal_name "yxn_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_39;// synopsys keep_signal_name "yxn_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_40;// synopsys keep_signal_name "yxn_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_41;// synopsys keep_signal_name "yxn_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_42;// synopsys keep_signal_name "yxn_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_43;// synopsys keep_signal_name "yxn_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_44;// synopsys keep_signal_name "yxn_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_45;// synopsys keep_signal_name "yxn_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_46;// synopsys keep_signal_name "yxn_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_47;// synopsys keep_signal_name "yxn_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_48;// synopsys keep_signal_name "yxn_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_49;// synopsys keep_signal_name "yxn_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_50;// synopsys keep_signal_name "yxn_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_51;// synopsys keep_signal_name "yxn_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_52;// synopsys keep_signal_name "yxn_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_53;// synopsys keep_signal_name "yxn_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_54;// synopsys keep_signal_name "yxn_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] yxn_55;// synopsys keep_signal_name "yxn_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_0;// synopsys keep_signal_name "v_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_1;// synopsys keep_signal_name "v_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_2;// synopsys keep_signal_name "v_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_3;// synopsys keep_signal_name "v_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_4;// synopsys keep_signal_name "v_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_5;// synopsys keep_signal_name "v_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_6;// synopsys keep_signal_name "v_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_7;// synopsys keep_signal_name "v_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_8;// synopsys keep_signal_name "v_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_9;// synopsys keep_signal_name "v_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_10;// synopsys keep_signal_name "v_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_11;// synopsys keep_signal_name "v_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_12;// synopsys keep_signal_name "v_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_13;// synopsys keep_signal_name "v_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_14;// synopsys keep_signal_name "v_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_15;// synopsys keep_signal_name "v_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_16;// synopsys keep_signal_name "v_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_17;// synopsys keep_signal_name "v_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_18;// synopsys keep_signal_name "v_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_19;// synopsys keep_signal_name "v_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_20;// synopsys keep_signal_name "v_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_21;// synopsys keep_signal_name "v_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_22;// synopsys keep_signal_name "v_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_23;// synopsys keep_signal_name "v_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_24;// synopsys keep_signal_name "v_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_25;// synopsys keep_signal_name "v_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_26;// synopsys keep_signal_name "v_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_27;// synopsys keep_signal_name "v_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_28;// synopsys keep_signal_name "v_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_29;// synopsys keep_signal_name "v_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_30;// synopsys keep_signal_name "v_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_31;// synopsys keep_signal_name "v_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_32;// synopsys keep_signal_name "v_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_33;// synopsys keep_signal_name "v_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_34;// synopsys keep_signal_name "v_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_35;// synopsys keep_signal_name "v_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_36;// synopsys keep_signal_name "v_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_37;// synopsys keep_signal_name "v_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_38;// synopsys keep_signal_name "v_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_39;// synopsys keep_signal_name "v_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_40;// synopsys keep_signal_name "v_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_41;// synopsys keep_signal_name "v_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_42;// synopsys keep_signal_name "v_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_43;// synopsys keep_signal_name "v_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_44;// synopsys keep_signal_name "v_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_45;// synopsys keep_signal_name "v_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_46;// synopsys keep_signal_name "v_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_47;// synopsys keep_signal_name "v_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_48;// synopsys keep_signal_name "v_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_49;// synopsys keep_signal_name "v_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_50;// synopsys keep_signal_name "v_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_51;// synopsys keep_signal_name "v_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_52;// synopsys keep_signal_name "v_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_53;// synopsys keep_signal_name "v_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_54;// synopsys keep_signal_name "v_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] v_55;// synopsys keep_signal_name "v_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire vldd2;
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_0;// synopsys keep_signal_name "xdn_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_1;// synopsys keep_signal_name "xdn_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_2;// synopsys keep_signal_name "xdn_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_3;// synopsys keep_signal_name "xdn_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_4;// synopsys keep_signal_name "xdn_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_5;// synopsys keep_signal_name "xdn_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_6;// synopsys keep_signal_name "xdn_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_7;// synopsys keep_signal_name "xdn_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_8;// synopsys keep_signal_name "xdn_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_9;// synopsys keep_signal_name "xdn_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_10;// synopsys keep_signal_name "xdn_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_11;// synopsys keep_signal_name "xdn_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_12;// synopsys keep_signal_name "xdn_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_13;// synopsys keep_signal_name "xdn_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_14;// synopsys keep_signal_name "xdn_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_15;// synopsys keep_signal_name "xdn_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_16;// synopsys keep_signal_name "xdn_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_17;// synopsys keep_signal_name "xdn_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_18;// synopsys keep_signal_name "xdn_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_19;// synopsys keep_signal_name "xdn_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_20;// synopsys keep_signal_name "xdn_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_21;// synopsys keep_signal_name "xdn_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_22;// synopsys keep_signal_name "xdn_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_23;// synopsys keep_signal_name "xdn_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_24;// synopsys keep_signal_name "xdn_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_25;// synopsys keep_signal_name "xdn_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_26;// synopsys keep_signal_name "xdn_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_27;// synopsys keep_signal_name "xdn_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_28;// synopsys keep_signal_name "xdn_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_29;// synopsys keep_signal_name "xdn_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_30;// synopsys keep_signal_name "xdn_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_31;// synopsys keep_signal_name "xdn_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_32;// synopsys keep_signal_name "xdn_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_33;// synopsys keep_signal_name "xdn_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_34;// synopsys keep_signal_name "xdn_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_35;// synopsys keep_signal_name "xdn_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_36;// synopsys keep_signal_name "xdn_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_37;// synopsys keep_signal_name "xdn_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_38;// synopsys keep_signal_name "xdn_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_39;// synopsys keep_signal_name "xdn_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_40;// synopsys keep_signal_name "xdn_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_41;// synopsys keep_signal_name "xdn_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_42;// synopsys keep_signal_name "xdn_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_43;// synopsys keep_signal_name "xdn_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_44;// synopsys keep_signal_name "xdn_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_45;// synopsys keep_signal_name "xdn_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_46;// synopsys keep_signal_name "xdn_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_47;// synopsys keep_signal_name "xdn_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_48;// synopsys keep_signal_name "xdn_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_49;// synopsys keep_signal_name "xdn_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_50;// synopsys keep_signal_name "xdn_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_51;// synopsys keep_signal_name "xdn_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_52;// synopsys keep_signal_name "xdn_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_53;// synopsys keep_signal_name "xdn_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_54;// synopsys keep_signal_name "xdn_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xdn_55;// synopsys keep_signal_name "xdn_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_0;// synopsys keep_signal_name "xar_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_1;// synopsys keep_signal_name "xar_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_2;// synopsys keep_signal_name "xar_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_3;// synopsys keep_signal_name "xar_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_4;// synopsys keep_signal_name "xar_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_5;// synopsys keep_signal_name "xar_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_6;// synopsys keep_signal_name "xar_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_7;// synopsys keep_signal_name "xar_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_8;// synopsys keep_signal_name "xar_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_9;// synopsys keep_signal_name "xar_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_10;// synopsys keep_signal_name "xar_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_11;// synopsys keep_signal_name "xar_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_12;// synopsys keep_signal_name "xar_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_13;// synopsys keep_signal_name "xar_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_14;// synopsys keep_signal_name "xar_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_15;// synopsys keep_signal_name "xar_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_16;// synopsys keep_signal_name "xar_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_17;// synopsys keep_signal_name "xar_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_18;// synopsys keep_signal_name "xar_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_19;// synopsys keep_signal_name "xar_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_20;// synopsys keep_signal_name "xar_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_21;// synopsys keep_signal_name "xar_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_22;// synopsys keep_signal_name "xar_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_23;// synopsys keep_signal_name "xar_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_24;// synopsys keep_signal_name "xar_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_25;// synopsys keep_signal_name "xar_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_26;// synopsys keep_signal_name "xar_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_27;// synopsys keep_signal_name "xar_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_28;// synopsys keep_signal_name "xar_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_29;// synopsys keep_signal_name "xar_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_30;// synopsys keep_signal_name "xar_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_31;// synopsys keep_signal_name "xar_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_32;// synopsys keep_signal_name "xar_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_33;// synopsys keep_signal_name "xar_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_34;// synopsys keep_signal_name "xar_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_35;// synopsys keep_signal_name "xar_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_36;// synopsys keep_signal_name "xar_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_37;// synopsys keep_signal_name "xar_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_38;// synopsys keep_signal_name "xar_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_39;// synopsys keep_signal_name "xar_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_40;// synopsys keep_signal_name "xar_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_41;// synopsys keep_signal_name "xar_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_42;// synopsys keep_signal_name "xar_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_43;// synopsys keep_signal_name "xar_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_44;// synopsys keep_signal_name "xar_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_45;// synopsys keep_signal_name "xar_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_46;// synopsys keep_signal_name "xar_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_47;// synopsys keep_signal_name "xar_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_48;// synopsys keep_signal_name "xar_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_49;// synopsys keep_signal_name "xar_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_50;// synopsys keep_signal_name "xar_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_51;// synopsys keep_signal_name "xar_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_52;// synopsys keep_signal_name "xar_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_53;// synopsys keep_signal_name "xar_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_54;// synopsys keep_signal_name "xar_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xar_55;// synopsys keep_signal_name "xar_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_0;// synopsys keep_signal_name "u_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_1;// synopsys keep_signal_name "u_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_2;// synopsys keep_signal_name "u_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_3;// synopsys keep_signal_name "u_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_4;// synopsys keep_signal_name "u_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_5;// synopsys keep_signal_name "u_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_6;// synopsys keep_signal_name "u_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_7;// synopsys keep_signal_name "u_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_8;// synopsys keep_signal_name "u_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_9;// synopsys keep_signal_name "u_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_10;// synopsys keep_signal_name "u_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_11;// synopsys keep_signal_name "u_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_12;// synopsys keep_signal_name "u_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_13;// synopsys keep_signal_name "u_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_14;// synopsys keep_signal_name "u_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_15;// synopsys keep_signal_name "u_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_16;// synopsys keep_signal_name "u_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_17;// synopsys keep_signal_name "u_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_18;// synopsys keep_signal_name "u_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_19;// synopsys keep_signal_name "u_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_20;// synopsys keep_signal_name "u_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_21;// synopsys keep_signal_name "u_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_22;// synopsys keep_signal_name "u_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_23;// synopsys keep_signal_name "u_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_24;// synopsys keep_signal_name "u_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_25;// synopsys keep_signal_name "u_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_26;// synopsys keep_signal_name "u_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_27;// synopsys keep_signal_name "u_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_28;// synopsys keep_signal_name "u_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_29;// synopsys keep_signal_name "u_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_30;// synopsys keep_signal_name "u_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_31;// synopsys keep_signal_name "u_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_32;// synopsys keep_signal_name "u_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_33;// synopsys keep_signal_name "u_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_34;// synopsys keep_signal_name "u_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_35;// synopsys keep_signal_name "u_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_36;// synopsys keep_signal_name "u_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_37;// synopsys keep_signal_name "u_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_38;// synopsys keep_signal_name "u_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_39;// synopsys keep_signal_name "u_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_40;// synopsys keep_signal_name "u_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_41;// synopsys keep_signal_name "u_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_42;// synopsys keep_signal_name "u_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_43;// synopsys keep_signal_name "u_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_44;// synopsys keep_signal_name "u_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_45;// synopsys keep_signal_name "u_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_46;// synopsys keep_signal_name "u_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_47;// synopsys keep_signal_name "u_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_48;// synopsys keep_signal_name "u_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_49;// synopsys keep_signal_name "u_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_50;// synopsys keep_signal_name "u_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_51;// synopsys keep_signal_name "u_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_52;// synopsys keep_signal_name "u_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_53;// synopsys keep_signal_name "u_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_54;// synopsys keep_signal_name "u_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] u_55;// synopsys keep_signal_name "u_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_0;// synopsys keep_signal_name "xay_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_1;// synopsys keep_signal_name "xay_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_2;// synopsys keep_signal_name "xay_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_3;// synopsys keep_signal_name "xay_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_4;// synopsys keep_signal_name "xay_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_5;// synopsys keep_signal_name "xay_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_6;// synopsys keep_signal_name "xay_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xay_7;// synopsys keep_signal_name "xay_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_0;// synopsys keep_signal_name "k_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_1;// synopsys keep_signal_name "k_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_2;// synopsys keep_signal_name "k_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_3;// synopsys keep_signal_name "k_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_4;// synopsys keep_signal_name "k_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_5;// synopsys keep_signal_name "k_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_6;// synopsys keep_signal_name "k_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] k_7;// synopsys keep_signal_name "k_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_0;// synopsys keep_signal_name "xav_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_1;// synopsys keep_signal_name "xav_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_2;// synopsys keep_signal_name "xav_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_3;// synopsys keep_signal_name "xav_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_4;// synopsys keep_signal_name "xav_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_5;// synopsys keep_signal_name "xav_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_6;// synopsys keep_signal_name "xav_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_7;// synopsys keep_signal_name "xav_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_8;// synopsys keep_signal_name "xav_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_9;// synopsys keep_signal_name "xav_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_10;// synopsys keep_signal_name "xav_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_11;// synopsys keep_signal_name "xav_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_12;// synopsys keep_signal_name "xav_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_13;// synopsys keep_signal_name "xav_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_14;// synopsys keep_signal_name "xav_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_15;// synopsys keep_signal_name "xav_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_16;// synopsys keep_signal_name "xav_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_17;// synopsys keep_signal_name "xav_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_18;// synopsys keep_signal_name "xav_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_19;// synopsys keep_signal_name "xav_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_20;// synopsys keep_signal_name "xav_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_21;// synopsys keep_signal_name "xav_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_22;// synopsys keep_signal_name "xav_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_23;// synopsys keep_signal_name "xav_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_24;// synopsys keep_signal_name "xav_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_25;// synopsys keep_signal_name "xav_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_26;// synopsys keep_signal_name "xav_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_27;// synopsys keep_signal_name "xav_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_28;// synopsys keep_signal_name "xav_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_29;// synopsys keep_signal_name "xav_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_30;// synopsys keep_signal_name "xav_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_31;// synopsys keep_signal_name "xav_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_32;// synopsys keep_signal_name "xav_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_33;// synopsys keep_signal_name "xav_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_34;// synopsys keep_signal_name "xav_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_35;// synopsys keep_signal_name "xav_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_36;// synopsys keep_signal_name "xav_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_37;// synopsys keep_signal_name "xav_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_38;// synopsys keep_signal_name "xav_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_39;// synopsys keep_signal_name "xav_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_40;// synopsys keep_signal_name "xav_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_41;// synopsys keep_signal_name "xav_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_42;// synopsys keep_signal_name "xav_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_43;// synopsys keep_signal_name "xav_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_44;// synopsys keep_signal_name "xav_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_45;// synopsys keep_signal_name "xav_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_46;// synopsys keep_signal_name "xav_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_47;// synopsys keep_signal_name "xav_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_48;// synopsys keep_signal_name "xav_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_49;// synopsys keep_signal_name "xav_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_50;// synopsys keep_signal_name "xav_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_51;// synopsys keep_signal_name "xav_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_52;// synopsys keep_signal_name "xav_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_53;// synopsys keep_signal_name "xav_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_54;// synopsys keep_signal_name "xav_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] xav_55;// synopsys keep_signal_name "xav_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_0;// synopsys keep_signal_name "t_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_1;// synopsys keep_signal_name "t_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_2;// synopsys keep_signal_name "t_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_3;// synopsys keep_signal_name "t_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_4;// synopsys keep_signal_name "t_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_5;// synopsys keep_signal_name "t_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_6;// synopsys keep_signal_name "t_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_7;// synopsys keep_signal_name "t_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_8;// synopsys keep_signal_name "t_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_9;// synopsys keep_signal_name "t_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_10;// synopsys keep_signal_name "t_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_11;// synopsys keep_signal_name "t_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_12;// synopsys keep_signal_name "t_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_13;// synopsys keep_signal_name "t_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_14;// synopsys keep_signal_name "t_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_15;// synopsys keep_signal_name "t_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_16;// synopsys keep_signal_name "t_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_17;// synopsys keep_signal_name "t_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_18;// synopsys keep_signal_name "t_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_19;// synopsys keep_signal_name "t_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_20;// synopsys keep_signal_name "t_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_21;// synopsys keep_signal_name "t_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_22;// synopsys keep_signal_name "t_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_23;// synopsys keep_signal_name "t_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_24;// synopsys keep_signal_name "t_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_25;// synopsys keep_signal_name "t_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_26;// synopsys keep_signal_name "t_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_27;// synopsys keep_signal_name "t_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_28;// synopsys keep_signal_name "t_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_29;// synopsys keep_signal_name "t_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_30;// synopsys keep_signal_name "t_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_31;// synopsys keep_signal_name "t_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_32;// synopsys keep_signal_name "t_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_33;// synopsys keep_signal_name "t_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_34;// synopsys keep_signal_name "t_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_35;// synopsys keep_signal_name "t_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_36;// synopsys keep_signal_name "t_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_37;// synopsys keep_signal_name "t_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_38;// synopsys keep_signal_name "t_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_39;// synopsys keep_signal_name "t_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_40;// synopsys keep_signal_name "t_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_41;// synopsys keep_signal_name "t_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_42;// synopsys keep_signal_name "t_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_43;// synopsys keep_signal_name "t_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_44;// synopsys keep_signal_name "t_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_45;// synopsys keep_signal_name "t_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_46;// synopsys keep_signal_name "t_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_47;// synopsys keep_signal_name "t_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_48;// synopsys keep_signal_name "t_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_49;// synopsys keep_signal_name "t_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_50;// synopsys keep_signal_name "t_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_51;// synopsys keep_signal_name "t_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_52;// synopsys keep_signal_name "t_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_53;// synopsys keep_signal_name "t_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_54;// synopsys keep_signal_name "t_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] t_55;// synopsys keep_signal_name "t_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_0;// synopsys keep_signal_name "z_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_1;// synopsys keep_signal_name "z_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_2;// synopsys keep_signal_name "z_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_3;// synopsys keep_signal_name "z_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_4;// synopsys keep_signal_name "z_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_5;// synopsys keep_signal_name "z_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_6;// synopsys keep_signal_name "z_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_7;// synopsys keep_signal_name "z_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_8;// synopsys keep_signal_name "z_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_9;// synopsys keep_signal_name "z_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_10;// synopsys keep_signal_name "z_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_11;// synopsys keep_signal_name "z_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_12;// synopsys keep_signal_name "z_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_13;// synopsys keep_signal_name "z_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_14;// synopsys keep_signal_name "z_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_15;// synopsys keep_signal_name "z_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_16;// synopsys keep_signal_name "z_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_17;// synopsys keep_signal_name "z_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_18;// synopsys keep_signal_name "z_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_19;// synopsys keep_signal_name "z_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_20;// synopsys keep_signal_name "z_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_21;// synopsys keep_signal_name "z_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_22;// synopsys keep_signal_name "z_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_23;// synopsys keep_signal_name "z_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_24;// synopsys keep_signal_name "z_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_25;// synopsys keep_signal_name "z_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_26;// synopsys keep_signal_name "z_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_27;// synopsys keep_signal_name "z_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_28;// synopsys keep_signal_name "z_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_29;// synopsys keep_signal_name "z_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_30;// synopsys keep_signal_name "z_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_31;// synopsys keep_signal_name "z_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_32;// synopsys keep_signal_name "z_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_33;// synopsys keep_signal_name "z_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_34;// synopsys keep_signal_name "z_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_35;// synopsys keep_signal_name "z_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_36;// synopsys keep_signal_name "z_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_37;// synopsys keep_signal_name "z_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_38;// synopsys keep_signal_name "z_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_39;// synopsys keep_signal_name "z_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_40;// synopsys keep_signal_name "z_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_41;// synopsys keep_signal_name "z_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_42;// synopsys keep_signal_name "z_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_43;// synopsys keep_signal_name "z_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_44;// synopsys keep_signal_name "z_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_45;// synopsys keep_signal_name "z_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_46;// synopsys keep_signal_name "z_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_47;// synopsys keep_signal_name "z_47"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_48;// synopsys keep_signal_name "z_48"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_49;// synopsys keep_signal_name "z_49"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_50;// synopsys keep_signal_name "z_50"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_51;// synopsys keep_signal_name "z_51"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_52;// synopsys keep_signal_name "z_52"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_53;// synopsys keep_signal_name "z_53"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_54;// synopsys keep_signal_name "z_54"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] z_55;// synopsys keep_signal_name "z_55"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_0;// synopsys keep_signal_name "zxz_0"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_1;// synopsys keep_signal_name "zxz_1"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_2;// synopsys keep_signal_name "zxz_2"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_3;// synopsys keep_signal_name "zxz_3"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_4;// synopsys keep_signal_name "zxz_4"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_5;// synopsys keep_signal_name "zxz_5"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_6;// synopsys keep_signal_name "zxz_6"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_7;// synopsys keep_signal_name "zxz_7"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_8;// synopsys keep_signal_name "zxz_8"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_9;// synopsys keep_signal_name "zxz_9"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_10;// synopsys keep_signal_name "zxz_10"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_11;// synopsys keep_signal_name "zxz_11"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_12;// synopsys keep_signal_name "zxz_12"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_13;// synopsys keep_signal_name "zxz_13"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_14;// synopsys keep_signal_name "zxz_14"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_15;// synopsys keep_signal_name "zxz_15"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_16;// synopsys keep_signal_name "zxz_16"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_17;// synopsys keep_signal_name "zxz_17"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_18;// synopsys keep_signal_name "zxz_18"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_19;// synopsys keep_signal_name "zxz_19"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_20;// synopsys keep_signal_name "zxz_20"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_21;// synopsys keep_signal_name "zxz_21"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_22;// synopsys keep_signal_name "zxz_22"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_23;// synopsys keep_signal_name "zxz_23"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_24;// synopsys keep_signal_name "zxz_24"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_25;// synopsys keep_signal_name "zxz_25"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_26;// synopsys keep_signal_name "zxz_26"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_27;// synopsys keep_signal_name "zxz_27"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_28;// synopsys keep_signal_name "zxz_28"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_29;// synopsys keep_signal_name "zxz_29"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_30;// synopsys keep_signal_name "zxz_30"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_31;// synopsys keep_signal_name "zxz_31"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_32;// synopsys keep_signal_name "zxz_32"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_33;// synopsys keep_signal_name "zxz_33"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_34;// synopsys keep_signal_name "zxz_34"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_35;// synopsys keep_signal_name "zxz_35"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_36;// synopsys keep_signal_name "zxz_36"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_37;// synopsys keep_signal_name "zxz_37"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_38;// synopsys keep_signal_name "zxz_38"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_39;// synopsys keep_signal_name "zxz_39"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_40;// synopsys keep_signal_name "zxz_40"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_41;// synopsys keep_signal_name "zxz_41"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_42;// synopsys keep_signal_name "zxz_42"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_43;// synopsys keep_signal_name "zxz_43"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_44;// synopsys keep_signal_name "zxz_44"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_45;// synopsys keep_signal_name "zxz_45"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_46;// synopsys keep_signal_name "zxz_46"
(*DONT_TOUCH="YES"*)(*KEEP="TRUE"*)wire [31:0] zxz_47;// synopsys keep_signal_name "zxz_47"

// delay i_dvld
lix_reg
  #(.W (1))
  u0_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (1'd1),
    .i_en   (i_rvld),
    .i_x    (i_dvld),
    .o_z    (vldd1));



// delay i_x[0+:32]
lix_reg
  #(.W (32))
  u1_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[0+:32]),
    .o_z    (xd_0));



// delay i_x[32+:32]
lix_reg
  #(.W (32))
  u2_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[32+:32]),
    .o_z    (xd_1));



// delay i_x[64+:32]
lix_reg
  #(.W (32))
  u3_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[64+:32]),
    .o_z    (xd_2));



// delay i_x[96+:32]
lix_reg
  #(.W (32))
  u4_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[96+:32]),
    .o_z    (xd_3));



// delay i_x[128+:32]
lix_reg
  #(.W (32))
  u5_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[128+:32]),
    .o_z    (xd_4));



// delay i_x[160+:32]
lix_reg
  #(.W (32))
  u6_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[160+:32]),
    .o_z    (xd_5));



// delay i_x[192+:32]
lix_reg
  #(.W (32))
  u7_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[192+:32]),
    .o_z    (xd_6));



// delay i_x[224+:32]
lix_reg
  #(.W (32))
  u8_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_x[224+:32]),
    .o_z    (xd_7));



// delay i_y[0+:32]
lix_reg
  #(.W (32))
  u9_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[0+:32]),
    .o_z    (yd_0));



// delay i_y[32+:32]
lix_reg
  #(.W (32))
  u10_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[32+:32]),
    .o_z    (yd_1));



// delay i_y[64+:32]
lix_reg
  #(.W (32))
  u11_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[64+:32]),
    .o_z    (yd_2));



// delay i_y[96+:32]
lix_reg
  #(.W (32))
  u12_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[96+:32]),
    .o_z    (yd_3));



// delay i_y[128+:32]
lix_reg
  #(.W (32))
  u13_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[128+:32]),
    .o_z    (yd_4));



// delay i_y[160+:32]
lix_reg
  #(.W (32))
  u14_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[160+:32]),
    .o_z    (yd_5));



// delay i_y[192+:32]
lix_reg
  #(.W (32))
  u15_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[192+:32]),
    .o_z    (yd_6));



// delay i_y[224+:32]
lix_reg
  #(.W (32))
  u16_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_y[224+:32]),
    .o_z    (yd_7));



// delay i_n0
lix_reg
  #(.W (32))
  u17_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[0+:32]),
    .o_z    (r_0));



// delay i_n1
lix_reg
  #(.W (32))
  u18_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[32+:32]),
    .o_z    (r_1));



// delay i_n2
lix_reg
  #(.W (32))
  u19_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[64+:32]),
    .o_z    (r_2));



// delay i_n3
lix_reg
  #(.W (32))
  u20_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[96+:32]),
    .o_z    (r_3));



// delay i_n4
lix_reg
  #(.W (32))
  u21_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[128+:32]),
    .o_z    (r_4));



// delay i_n5
lix_reg
  #(.W (32))
  u22_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[160+:32]),
    .o_z    (r_5));



// delay i_n6
lix_reg
  #(.W (32))
  u23_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[192+:32]),
    .o_z    (r_6));



// delay i_n0
lix_reg
  #(.W (32))
  u24_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[0+:32]),
    .o_z    (r_7));



// delay i_n7
lix_reg
  #(.W (32))
  u25_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[224+:32]),
    .o_z    (r_8));



// delay i_n8
lix_reg
  #(.W (32))
  u26_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[256+:32]),
    .o_z    (r_9));



// delay i_n9
lix_reg
  #(.W (32))
  u27_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[288+:32]),
    .o_z    (r_10));



// delay i_n10
lix_reg
  #(.W (32))
  u28_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[320+:32]),
    .o_z    (r_11));



// delay i_n11
lix_reg
  #(.W (32))
  u29_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[352+:32]),
    .o_z    (r_12));



// delay i_n12
lix_reg
  #(.W (32))
  u30_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[384+:32]),
    .o_z    (r_13));



// delay i_n1
lix_reg
  #(.W (32))
  u31_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[32+:32]),
    .o_z    (r_14));



// delay i_n7
lix_reg
  #(.W (32))
  u32_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[224+:32]),
    .o_z    (r_15));



// delay i_n13
lix_reg
  #(.W (32))
  u33_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[416+:32]),
    .o_z    (r_16));



// delay i_n14
lix_reg
  #(.W (32))
  u34_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[448+:32]),
    .o_z    (r_17));



// delay i_n15
lix_reg
  #(.W (32))
  u35_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[480+:32]),
    .o_z    (r_18));



// delay i_n16
lix_reg
  #(.W (32))
  u36_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[512+:32]),
    .o_z    (r_19));



// delay i_n17
lix_reg
  #(.W (32))
  u37_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[544+:32]),
    .o_z    (r_20));



// delay i_n2
lix_reg
  #(.W (32))
  u38_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[64+:32]),
    .o_z    (r_21));



// delay i_n8
lix_reg
  #(.W (32))
  u39_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[256+:32]),
    .o_z    (r_22));



// delay i_n13
lix_reg
  #(.W (32))
  u40_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[416+:32]),
    .o_z    (r_23));



// delay i_n18
lix_reg
  #(.W (32))
  u41_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[576+:32]),
    .o_z    (r_24));



// delay i_n19
lix_reg
  #(.W (32))
  u42_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[608+:32]),
    .o_z    (r_25));



// delay i_n20
lix_reg
  #(.W (32))
  u43_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[640+:32]),
    .o_z    (r_26));



// delay i_n21
lix_reg
  #(.W (32))
  u44_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[672+:32]),
    .o_z    (r_27));



// delay i_n3
lix_reg
  #(.W (32))
  u45_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[96+:32]),
    .o_z    (r_28));



// delay i_n9
lix_reg
  #(.W (32))
  u46_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[288+:32]),
    .o_z    (r_29));



// delay i_n14
lix_reg
  #(.W (32))
  u47_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[448+:32]),
    .o_z    (r_30));



// delay i_n18
lix_reg
  #(.W (32))
  u48_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[576+:32]),
    .o_z    (r_31));



// delay i_n22
lix_reg
  #(.W (32))
  u49_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[704+:32]),
    .o_z    (r_32));



// delay i_n23
lix_reg
  #(.W (32))
  u50_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[736+:32]),
    .o_z    (r_33));



// delay i_n24
lix_reg
  #(.W (32))
  u51_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[768+:32]),
    .o_z    (r_34));



// delay i_n4
lix_reg
  #(.W (32))
  u52_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[128+:32]),
    .o_z    (r_35));



// delay i_n10
lix_reg
  #(.W (32))
  u53_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[320+:32]),
    .o_z    (r_36));



// delay i_n15
lix_reg
  #(.W (32))
  u54_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[480+:32]),
    .o_z    (r_37));



// delay i_n19
lix_reg
  #(.W (32))
  u55_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[608+:32]),
    .o_z    (r_38));



// delay i_n22
lix_reg
  #(.W (32))
  u56_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[704+:32]),
    .o_z    (r_39));



// delay i_n25
lix_reg
  #(.W (32))
  u57_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[800+:32]),
    .o_z    (r_40));



// delay i_n26
lix_reg
  #(.W (32))
  u58_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[832+:32]),
    .o_z    (r_41));



// delay i_n5
lix_reg
  #(.W (32))
  u59_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[160+:32]),
    .o_z    (r_42));



// delay i_n11
lix_reg
  #(.W (32))
  u60_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[352+:32]),
    .o_z    (r_43));



// delay i_n16
lix_reg
  #(.W (32))
  u61_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[512+:32]),
    .o_z    (r_44));



// delay i_n20
lix_reg
  #(.W (32))
  u62_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[640+:32]),
    .o_z    (r_45));



// delay i_n23
lix_reg
  #(.W (32))
  u63_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[736+:32]),
    .o_z    (r_46));



// delay i_n25
lix_reg
  #(.W (32))
  u64_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[800+:32]),
    .o_z    (r_47));



// delay i_n27
lix_reg
  #(.W (32))
  u65_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[864+:32]),
    .o_z    (r_48));



// delay i_n6
lix_reg
  #(.W (32))
  u66_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[192+:32]),
    .o_z    (r_49));



// delay i_n12
lix_reg
  #(.W (32))
  u67_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[384+:32]),
    .o_z    (r_50));



// delay i_n17
lix_reg
  #(.W (32))
  u68_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[544+:32]),
    .o_z    (r_51));



// delay i_n21
lix_reg
  #(.W (32))
  u69_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[672+:32]),
    .o_z    (r_52));



// delay i_n24
lix_reg
  #(.W (32))
  u70_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[768+:32]),
    .o_z    (r_53));



// delay i_n26
lix_reg
  #(.W (32))
  u71_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[832+:32]),
    .o_z    (r_54));



// delay i_n27
lix_reg
  #(.W (32))
  u72_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (i_n[864+:32]),
    .o_z    (r_55));



// i_y[0+:32] ^ i_n[0+:32]
lix_xor
  #(.W (32))
  u73_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[0+:32]),
    .o_z (yxn_0));



// i_y[0+:32] ^ i_n[32+:32]
lix_xor
  #(.W (32))
  u74_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[32+:32]),
    .o_z (yxn_1));



// i_y[0+:32] ^ i_n[64+:32]
lix_xor
  #(.W (32))
  u75_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[64+:32]),
    .o_z (yxn_2));



// i_y[0+:32] ^ i_n[96+:32]
lix_xor
  #(.W (32))
  u76_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[96+:32]),
    .o_z (yxn_3));



// i_y[0+:32] ^ i_n[128+:32]
lix_xor
  #(.W (32))
  u77_lix_xor
   (.i_x (i_y[160+:32]),
    .i_y (i_n[128+:32]),
    .o_z (yxn_4));



// i_y[0+:32] ^ i_n[160+:32]
lix_xor
  #(.W (32))
  u78_lix_xor
   (.i_x (i_y[192+:32]),
    .i_y (i_n[160+:32]),
    .o_z (yxn_5));



// i_y[0+:32] ^ i_n[192+:32]
lix_xor
  #(.W (32))
  u79_lix_xor
   (.i_x (i_y[224+:32]),
    .i_y (i_n[192+:32]),
    .o_z (yxn_6));



// i_y[32+:32] ^ i_n[0+:32]
lix_xor
  #(.W (32))
  u80_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[0+:32]),
    .o_z (yxn_7));



// i_y[32+:32] ^ i_n[224+:32]
lix_xor
  #(.W (32))
  u81_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[224+:32]),
    .o_z (yxn_8));



// i_y[32+:32] ^ i_n[256+:32]
lix_xor
  #(.W (32))
  u82_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[256+:32]),
    .o_z (yxn_9));



// i_y[32+:32] ^ i_n[288+:32]
lix_xor
  #(.W (32))
  u83_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[288+:32]),
    .o_z (yxn_10));



// i_y[32+:32] ^ i_n[320+:32]
lix_xor
  #(.W (32))
  u84_lix_xor
   (.i_x (i_y[160+:32]),
    .i_y (i_n[320+:32]),
    .o_z (yxn_11));



// i_y[32+:32] ^ i_n[352+:32]
lix_xor
  #(.W (32))
  u85_lix_xor
   (.i_x (i_y[192+:32]),
    .i_y (i_n[352+:32]),
    .o_z (yxn_12));



// i_y[32+:32] ^ i_n[384+:32]
lix_xor
  #(.W (32))
  u86_lix_xor
   (.i_x (i_y[224+:32]),
    .i_y (i_n[384+:32]),
    .o_z (yxn_13));



// i_y[64+:32] ^ i_n[32+:32]
lix_xor
  #(.W (32))
  u87_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[32+:32]),
    .o_z (yxn_14));



// i_y[64+:32] ^ i_n[224+:32]
lix_xor
  #(.W (32))
  u88_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[224+:32]),
    .o_z (yxn_15));



// i_y[64+:32] ^ i_n[416+:32]
lix_xor
  #(.W (32))
  u89_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[416+:32]),
    .o_z (yxn_16));



// i_y[64+:32] ^ i_n[448+:32]
lix_xor
  #(.W (32))
  u90_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[448+:32]),
    .o_z (yxn_17));



// i_y[64+:32] ^ i_n[480+:32]
lix_xor
  #(.W (32))
  u91_lix_xor
   (.i_x (i_y[160+:32]),
    .i_y (i_n[480+:32]),
    .o_z (yxn_18));



// i_y[64+:32] ^ i_n[512+:32]
lix_xor
  #(.W (32))
  u92_lix_xor
   (.i_x (i_y[192+:32]),
    .i_y (i_n[512+:32]),
    .o_z (yxn_19));



// i_y[64+:32] ^ i_n[544+:32]
lix_xor
  #(.W (32))
  u93_lix_xor
   (.i_x (i_y[224+:32]),
    .i_y (i_n[544+:32]),
    .o_z (yxn_20));



// i_y[96+:32] ^ i_n[64+:32]
lix_xor
  #(.W (32))
  u94_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[64+:32]),
    .o_z (yxn_21));



// i_y[96+:32] ^ i_n[256+:32]
lix_xor
  #(.W (32))
  u95_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[256+:32]),
    .o_z (yxn_22));



// i_y[96+:32] ^ i_n[416+:32]
lix_xor
  #(.W (32))
  u96_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[416+:32]),
    .o_z (yxn_23));



// i_y[96+:32] ^ i_n[576+:32]
lix_xor
  #(.W (32))
  u97_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[576+:32]),
    .o_z (yxn_24));



// i_y[96+:32] ^ i_n[608+:32]
lix_xor
  #(.W (32))
  u98_lix_xor
   (.i_x (i_y[160+:32]),
    .i_y (i_n[608+:32]),
    .o_z (yxn_25));



// i_y[96+:32] ^ i_n[640+:32]
lix_xor
  #(.W (32))
  u99_lix_xor
   (.i_x (i_y[192+:32]),
    .i_y (i_n[640+:32]),
    .o_z (yxn_26));



// i_y[96+:32] ^ i_n[672+:32]
lix_xor
  #(.W (32))
  u100_lix_xor
   (.i_x (i_y[224+:32]),
    .i_y (i_n[672+:32]),
    .o_z (yxn_27));



// i_y[128+:32] ^ i_n[96+:32]
lix_xor
  #(.W (32))
  u101_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[96+:32]),
    .o_z (yxn_28));



// i_y[128+:32] ^ i_n[288+:32]
lix_xor
  #(.W (32))
  u102_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[288+:32]),
    .o_z (yxn_29));



// i_y[128+:32] ^ i_n[448+:32]
lix_xor
  #(.W (32))
  u103_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[448+:32]),
    .o_z (yxn_30));



// i_y[128+:32] ^ i_n[576+:32]
lix_xor
  #(.W (32))
  u104_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[576+:32]),
    .o_z (yxn_31));



// i_y[128+:32] ^ i_n[704+:32]
lix_xor
  #(.W (32))
  u105_lix_xor
   (.i_x (i_y[160+:32]),
    .i_y (i_n[704+:32]),
    .o_z (yxn_32));



// i_y[128+:32] ^ i_n[736+:32]
lix_xor
  #(.W (32))
  u106_lix_xor
   (.i_x (i_y[192+:32]),
    .i_y (i_n[736+:32]),
    .o_z (yxn_33));



// i_y[128+:32] ^ i_n[768+:32]
lix_xor
  #(.W (32))
  u107_lix_xor
   (.i_x (i_y[224+:32]),
    .i_y (i_n[768+:32]),
    .o_z (yxn_34));



// i_y[160+:32] ^ i_n[128+:32]
lix_xor
  #(.W (32))
  u108_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[128+:32]),
    .o_z (yxn_35));



// i_y[160+:32] ^ i_n[320+:32]
lix_xor
  #(.W (32))
  u109_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[320+:32]),
    .o_z (yxn_36));



// i_y[160+:32] ^ i_n[480+:32]
lix_xor
  #(.W (32))
  u110_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[480+:32]),
    .o_z (yxn_37));



// i_y[160+:32] ^ i_n[608+:32]
lix_xor
  #(.W (32))
  u111_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[608+:32]),
    .o_z (yxn_38));



// i_y[160+:32] ^ i_n[704+:32]
lix_xor
  #(.W (32))
  u112_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[704+:32]),
    .o_z (yxn_39));



// i_y[160+:32] ^ i_n[800+:32]
lix_xor
  #(.W (32))
  u113_lix_xor
   (.i_x (i_y[192+:32]),
    .i_y (i_n[800+:32]),
    .o_z (yxn_40));



// i_y[160+:32] ^ i_n[832+:32]
lix_xor
  #(.W (32))
  u114_lix_xor
   (.i_x (i_y[224+:32]),
    .i_y (i_n[832+:32]),
    .o_z (yxn_41));



// i_y[192+:32] ^ i_n[160+:32]
lix_xor
  #(.W (32))
  u115_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[160+:32]),
    .o_z (yxn_42));



// i_y[192+:32] ^ i_n[352+:32]
lix_xor
  #(.W (32))
  u116_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[352+:32]),
    .o_z (yxn_43));



// i_y[192+:32] ^ i_n[512+:32]
lix_xor
  #(.W (32))
  u117_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[512+:32]),
    .o_z (yxn_44));



// i_y[192+:32] ^ i_n[640+:32]
lix_xor
  #(.W (32))
  u118_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[640+:32]),
    .o_z (yxn_45));



// i_y[192+:32] ^ i_n[736+:32]
lix_xor
  #(.W (32))
  u119_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[736+:32]),
    .o_z (yxn_46));



// i_y[192+:32] ^ i_n[800+:32]
lix_xor
  #(.W (32))
  u120_lix_xor
   (.i_x (i_y[160+:32]),
    .i_y (i_n[800+:32]),
    .o_z (yxn_47));



// i_y[192+:32] ^ i_n[864+:32]
lix_xor
  #(.W (32))
  u121_lix_xor
   (.i_x (i_y[224+:32]),
    .i_y (i_n[864+:32]),
    .o_z (yxn_48));



// i_y[224+:32] ^ i_n[192+:32]
lix_xor
  #(.W (32))
  u122_lix_xor
   (.i_x (i_y[0+:32]),
    .i_y (i_n[192+:32]),
    .o_z (yxn_49));



// i_y[224+:32] ^ i_n[384+:32]
lix_xor
  #(.W (32))
  u123_lix_xor
   (.i_x (i_y[32+:32]),
    .i_y (i_n[384+:32]),
    .o_z (yxn_50));



// i_y[224+:32] ^ i_n[544+:32]
lix_xor
  #(.W (32))
  u124_lix_xor
   (.i_x (i_y[64+:32]),
    .i_y (i_n[544+:32]),
    .o_z (yxn_51));



// i_y[224+:32] ^ i_n[672+:32]
lix_xor
  #(.W (32))
  u125_lix_xor
   (.i_x (i_y[96+:32]),
    .i_y (i_n[672+:32]),
    .o_z (yxn_52));



// i_y[224+:32] ^ i_n[768+:32]
lix_xor
  #(.W (32))
  u126_lix_xor
   (.i_x (i_y[128+:32]),
    .i_y (i_n[768+:32]),
    .o_z (yxn_53));



// i_y[224+:32] ^ i_n[832+:32]
lix_xor
  #(.W (32))
  u127_lix_xor
   (.i_x (i_y[160+:32]),
    .i_y (i_n[832+:32]),
    .o_z (yxn_54));



// i_y[224+:32] ^ i_n[864+:32]
lix_xor
  #(.W (32))
  u128_lix_xor
   (.i_x (i_y[192+:32]),
    .i_y (i_n[864+:32]),
    .o_z (yxn_55));



// delay yxn_0
lix_reg
  #(.W (32))
  u129_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_0),
    .o_z    (v_0));



// delay yxn_1
lix_reg
  #(.W (32))
  u130_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_1),
    .o_z    (v_1));



// delay yxn_2
lix_reg
  #(.W (32))
  u131_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_2),
    .o_z    (v_2));



// delay yxn_3
lix_reg
  #(.W (32))
  u132_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_3),
    .o_z    (v_3));



// delay yxn_4
lix_reg
  #(.W (32))
  u133_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_4),
    .o_z    (v_4));



// delay yxn_5
lix_reg
  #(.W (32))
  u134_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_5),
    .o_z    (v_5));



// delay yxn_6
lix_reg
  #(.W (32))
  u135_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_6),
    .o_z    (v_6));



// delay yxn_7
lix_reg
  #(.W (32))
  u136_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_7),
    .o_z    (v_7));



// delay yxn_8
lix_reg
  #(.W (32))
  u137_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_8),
    .o_z    (v_8));



// delay yxn_9
lix_reg
  #(.W (32))
  u138_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_9),
    .o_z    (v_9));



// delay yxn_10
lix_reg
  #(.W (32))
  u139_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_10),
    .o_z    (v_10));



// delay yxn_11
lix_reg
  #(.W (32))
  u140_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_11),
    .o_z    (v_11));



// delay yxn_12
lix_reg
  #(.W (32))
  u141_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_12),
    .o_z    (v_12));



// delay yxn_13
lix_reg
  #(.W (32))
  u142_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_13),
    .o_z    (v_13));



// delay yxn_14
lix_reg
  #(.W (32))
  u143_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_14),
    .o_z    (v_14));



// delay yxn_15
lix_reg
  #(.W (32))
  u144_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_15),
    .o_z    (v_15));



// delay yxn_16
lix_reg
  #(.W (32))
  u145_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_16),
    .o_z    (v_16));



// delay yxn_17
lix_reg
  #(.W (32))
  u146_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_17),
    .o_z    (v_17));



// delay yxn_18
lix_reg
  #(.W (32))
  u147_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_18),
    .o_z    (v_18));



// delay yxn_19
lix_reg
  #(.W (32))
  u148_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_19),
    .o_z    (v_19));



// delay yxn_20
lix_reg
  #(.W (32))
  u149_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_20),
    .o_z    (v_20));



// delay yxn_21
lix_reg
  #(.W (32))
  u150_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_21),
    .o_z    (v_21));



// delay yxn_22
lix_reg
  #(.W (32))
  u151_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_22),
    .o_z    (v_22));



// delay yxn_23
lix_reg
  #(.W (32))
  u152_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_23),
    .o_z    (v_23));



// delay yxn_24
lix_reg
  #(.W (32))
  u153_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_24),
    .o_z    (v_24));



// delay yxn_25
lix_reg
  #(.W (32))
  u154_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_25),
    .o_z    (v_25));



// delay yxn_26
lix_reg
  #(.W (32))
  u155_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_26),
    .o_z    (v_26));



// delay yxn_27
lix_reg
  #(.W (32))
  u156_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_27),
    .o_z    (v_27));



// delay yxn_28
lix_reg
  #(.W (32))
  u157_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_28),
    .o_z    (v_28));



// delay yxn_29
lix_reg
  #(.W (32))
  u158_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_29),
    .o_z    (v_29));



// delay yxn_30
lix_reg
  #(.W (32))
  u159_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_30),
    .o_z    (v_30));



// delay yxn_31
lix_reg
  #(.W (32))
  u160_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_31),
    .o_z    (v_31));



// delay yxn_32
lix_reg
  #(.W (32))
  u161_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_32),
    .o_z    (v_32));



// delay yxn_33
lix_reg
  #(.W (32))
  u162_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_33),
    .o_z    (v_33));



// delay yxn_34
lix_reg
  #(.W (32))
  u163_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_34),
    .o_z    (v_34));



// delay yxn_35
lix_reg
  #(.W (32))
  u164_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_35),
    .o_z    (v_35));



// delay yxn_36
lix_reg
  #(.W (32))
  u165_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_36),
    .o_z    (v_36));



// delay yxn_37
lix_reg
  #(.W (32))
  u166_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_37),
    .o_z    (v_37));



// delay yxn_38
lix_reg
  #(.W (32))
  u167_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_38),
    .o_z    (v_38));



// delay yxn_39
lix_reg
  #(.W (32))
  u168_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_39),
    .o_z    (v_39));



// delay yxn_40
lix_reg
  #(.W (32))
  u169_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_40),
    .o_z    (v_40));



// delay yxn_41
lix_reg
  #(.W (32))
  u170_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_41),
    .o_z    (v_41));



// delay yxn_42
lix_reg
  #(.W (32))
  u171_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_42),
    .o_z    (v_42));



// delay yxn_43
lix_reg
  #(.W (32))
  u172_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_43),
    .o_z    (v_43));



// delay yxn_44
lix_reg
  #(.W (32))
  u173_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_44),
    .o_z    (v_44));



// delay yxn_45
lix_reg
  #(.W (32))
  u174_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_45),
    .o_z    (v_45));



// delay yxn_46
lix_reg
  #(.W (32))
  u175_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_46),
    .o_z    (v_46));



// delay yxn_47
lix_reg
  #(.W (32))
  u176_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_47),
    .o_z    (v_47));



// delay yxn_48
lix_reg
  #(.W (32))
  u177_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_48),
    .o_z    (v_48));



// delay yxn_49
lix_reg
  #(.W (32))
  u178_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_49),
    .o_z    (v_49));



// delay yxn_50
lix_reg
  #(.W (32))
  u179_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_50),
    .o_z    (v_50));



// delay yxn_51
lix_reg
  #(.W (32))
  u180_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_51),
    .o_z    (v_51));



// delay yxn_52
lix_reg
  #(.W (32))
  u181_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_52),
    .o_z    (v_52));



// delay yxn_53
lix_reg
  #(.W (32))
  u182_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_53),
    .o_z    (v_53));



// delay yxn_54
lix_reg
  #(.W (32))
  u183_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_54),
    .o_z    (v_54));



// delay yxn_55
lix_reg
  #(.W (32))
  u184_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (i_dvld),
    .i_en   (i_rvld),
    .i_x    (yxn_55),
    .o_z    (v_55));



// delay vldd1
lix_reg
  #(.W (1))
  u185_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (1'd1),
    .i_en   (i_rvld),
    .i_x    (vldd1),
    .o_z    (vldd2));



// not  xd_0
lix_not
  #(.W (32))
  u186_lix_not
   (.i_x (xd_0),
    .o_z (xdn_0));



// not  xd_1
lix_not
  #(.W (32))
  u187_lix_not
   (.i_x (xd_1),
    .o_z (xdn_1));



// not  xd_2
lix_not
  #(.W (32))
  u188_lix_not
   (.i_x (xd_2),
    .o_z (xdn_2));



// not  xd_3
lix_not
  #(.W (32))
  u189_lix_not
   (.i_x (xd_3),
    .o_z (xdn_3));



// not  xd_4
lix_not
  #(.W (32))
  u190_lix_not
   (.i_x (xd_4),
    .o_z (xdn_4));



// not  xd_5
lix_not
  #(.W (32))
  u191_lix_not
   (.i_x (xd_5),
    .o_z (xdn_5));



// not  xd_6
lix_not
  #(.W (32))
  u192_lix_not
   (.i_x (xd_6),
    .o_z (xdn_6));



// not  xd_7
lix_not
  #(.W (32))
  u193_lix_not
   (.i_x (xd_7),
    .o_z (xdn_7));



// ~xd_0 & r_0
lix_and
  #(.W (32))
  u194_lix_and
   (.i_x (xdn_0),
    .i_y (r_0),
    .o_z (xar_0));



// ~xd_0 & r_1
lix_and
  #(.W (32))
  u195_lix_and
   (.i_x (xdn_0),
    .i_y (r_1),
    .o_z (xar_1));



// ~xd_0 & r_2
lix_and
  #(.W (32))
  u196_lix_and
   (.i_x (xdn_0),
    .i_y (r_2),
    .o_z (xar_2));



// ~xd_0 & r_3
lix_and
  #(.W (32))
  u197_lix_and
   (.i_x (xdn_0),
    .i_y (r_3),
    .o_z (xar_3));



// ~xd_0 & r_4
lix_and
  #(.W (32))
  u198_lix_and
   (.i_x (xdn_0),
    .i_y (r_4),
    .o_z (xar_4));



// ~xd_0 & r_5
lix_and
  #(.W (32))
  u199_lix_and
   (.i_x (xdn_0),
    .i_y (r_5),
    .o_z (xar_5));



// ~xd_0 & r_6
lix_and
  #(.W (32))
  u200_lix_and
   (.i_x (xdn_0),
    .i_y (r_6),
    .o_z (xar_6));



// ~xd_1 & r_7
lix_and
  #(.W (32))
  u201_lix_and
   (.i_x (xdn_1),
    .i_y (r_7),
    .o_z (xar_7));



// ~xd_1 & r_8
lix_and
  #(.W (32))
  u202_lix_and
   (.i_x (xdn_1),
    .i_y (r_8),
    .o_z (xar_8));



// ~xd_1 & r_9
lix_and
  #(.W (32))
  u203_lix_and
   (.i_x (xdn_1),
    .i_y (r_9),
    .o_z (xar_9));



// ~xd_1 & r_10
lix_and
  #(.W (32))
  u204_lix_and
   (.i_x (xdn_1),
    .i_y (r_10),
    .o_z (xar_10));



// ~xd_1 & r_11
lix_and
  #(.W (32))
  u205_lix_and
   (.i_x (xdn_1),
    .i_y (r_11),
    .o_z (xar_11));



// ~xd_1 & r_12
lix_and
  #(.W (32))
  u206_lix_and
   (.i_x (xdn_1),
    .i_y (r_12),
    .o_z (xar_12));



// ~xd_1 & r_13
lix_and
  #(.W (32))
  u207_lix_and
   (.i_x (xdn_1),
    .i_y (r_13),
    .o_z (xar_13));



// ~xd_2 & r_14
lix_and
  #(.W (32))
  u208_lix_and
   (.i_x (xdn_2),
    .i_y (r_14),
    .o_z (xar_14));



// ~xd_2 & r_15
lix_and
  #(.W (32))
  u209_lix_and
   (.i_x (xdn_2),
    .i_y (r_15),
    .o_z (xar_15));



// ~xd_2 & r_16
lix_and
  #(.W (32))
  u210_lix_and
   (.i_x (xdn_2),
    .i_y (r_16),
    .o_z (xar_16));



// ~xd_2 & r_17
lix_and
  #(.W (32))
  u211_lix_and
   (.i_x (xdn_2),
    .i_y (r_17),
    .o_z (xar_17));



// ~xd_2 & r_18
lix_and
  #(.W (32))
  u212_lix_and
   (.i_x (xdn_2),
    .i_y (r_18),
    .o_z (xar_18));



// ~xd_2 & r_19
lix_and
  #(.W (32))
  u213_lix_and
   (.i_x (xdn_2),
    .i_y (r_19),
    .o_z (xar_19));



// ~xd_2 & r_20
lix_and
  #(.W (32))
  u214_lix_and
   (.i_x (xdn_2),
    .i_y (r_20),
    .o_z (xar_20));



// ~xd_3 & r_21
lix_and
  #(.W (32))
  u215_lix_and
   (.i_x (xdn_3),
    .i_y (r_21),
    .o_z (xar_21));



// ~xd_3 & r_22
lix_and
  #(.W (32))
  u216_lix_and
   (.i_x (xdn_3),
    .i_y (r_22),
    .o_z (xar_22));



// ~xd_3 & r_23
lix_and
  #(.W (32))
  u217_lix_and
   (.i_x (xdn_3),
    .i_y (r_23),
    .o_z (xar_23));



// ~xd_3 & r_24
lix_and
  #(.W (32))
  u218_lix_and
   (.i_x (xdn_3),
    .i_y (r_24),
    .o_z (xar_24));



// ~xd_3 & r_25
lix_and
  #(.W (32))
  u219_lix_and
   (.i_x (xdn_3),
    .i_y (r_25),
    .o_z (xar_25));



// ~xd_3 & r_26
lix_and
  #(.W (32))
  u220_lix_and
   (.i_x (xdn_3),
    .i_y (r_26),
    .o_z (xar_26));



// ~xd_3 & r_27
lix_and
  #(.W (32))
  u221_lix_and
   (.i_x (xdn_3),
    .i_y (r_27),
    .o_z (xar_27));



// ~xd_4 & r_28
lix_and
  #(.W (32))
  u222_lix_and
   (.i_x (xdn_4),
    .i_y (r_28),
    .o_z (xar_28));



// ~xd_4 & r_29
lix_and
  #(.W (32))
  u223_lix_and
   (.i_x (xdn_4),
    .i_y (r_29),
    .o_z (xar_29));



// ~xd_4 & r_30
lix_and
  #(.W (32))
  u224_lix_and
   (.i_x (xdn_4),
    .i_y (r_30),
    .o_z (xar_30));



// ~xd_4 & r_31
lix_and
  #(.W (32))
  u225_lix_and
   (.i_x (xdn_4),
    .i_y (r_31),
    .o_z (xar_31));



// ~xd_4 & r_32
lix_and
  #(.W (32))
  u226_lix_and
   (.i_x (xdn_4),
    .i_y (r_32),
    .o_z (xar_32));



// ~xd_4 & r_33
lix_and
  #(.W (32))
  u227_lix_and
   (.i_x (xdn_4),
    .i_y (r_33),
    .o_z (xar_33));



// ~xd_4 & r_34
lix_and
  #(.W (32))
  u228_lix_and
   (.i_x (xdn_4),
    .i_y (r_34),
    .o_z (xar_34));



// ~xd_5 & r_35
lix_and
  #(.W (32))
  u229_lix_and
   (.i_x (xdn_5),
    .i_y (r_35),
    .o_z (xar_35));



// ~xd_5 & r_36
lix_and
  #(.W (32))
  u230_lix_and
   (.i_x (xdn_5),
    .i_y (r_36),
    .o_z (xar_36));



// ~xd_5 & r_37
lix_and
  #(.W (32))
  u231_lix_and
   (.i_x (xdn_5),
    .i_y (r_37),
    .o_z (xar_37));



// ~xd_5 & r_38
lix_and
  #(.W (32))
  u232_lix_and
   (.i_x (xdn_5),
    .i_y (r_38),
    .o_z (xar_38));



// ~xd_5 & r_39
lix_and
  #(.W (32))
  u233_lix_and
   (.i_x (xdn_5),
    .i_y (r_39),
    .o_z (xar_39));



// ~xd_5 & r_40
lix_and
  #(.W (32))
  u234_lix_and
   (.i_x (xdn_5),
    .i_y (r_40),
    .o_z (xar_40));



// ~xd_5 & r_41
lix_and
  #(.W (32))
  u235_lix_and
   (.i_x (xdn_5),
    .i_y (r_41),
    .o_z (xar_41));



// ~xd_6 & r_42
lix_and
  #(.W (32))
  u236_lix_and
   (.i_x (xdn_6),
    .i_y (r_42),
    .o_z (xar_42));



// ~xd_6 & r_43
lix_and
  #(.W (32))
  u237_lix_and
   (.i_x (xdn_6),
    .i_y (r_43),
    .o_z (xar_43));



// ~xd_6 & r_44
lix_and
  #(.W (32))
  u238_lix_and
   (.i_x (xdn_6),
    .i_y (r_44),
    .o_z (xar_44));



// ~xd_6 & r_45
lix_and
  #(.W (32))
  u239_lix_and
   (.i_x (xdn_6),
    .i_y (r_45),
    .o_z (xar_45));



// ~xd_6 & r_46
lix_and
  #(.W (32))
  u240_lix_and
   (.i_x (xdn_6),
    .i_y (r_46),
    .o_z (xar_46));



// ~xd_6 & r_47
lix_and
  #(.W (32))
  u241_lix_and
   (.i_x (xdn_6),
    .i_y (r_47),
    .o_z (xar_47));



// ~xd_6 & r_48
lix_and
  #(.W (32))
  u242_lix_and
   (.i_x (xdn_6),
    .i_y (r_48),
    .o_z (xar_48));



// ~xd_7 & r_49
lix_and
  #(.W (32))
  u243_lix_and
   (.i_x (xdn_7),
    .i_y (r_49),
    .o_z (xar_49));



// ~xd_7 & r_50
lix_and
  #(.W (32))
  u244_lix_and
   (.i_x (xdn_7),
    .i_y (r_50),
    .o_z (xar_50));



// ~xd_7 & r_51
lix_and
  #(.W (32))
  u245_lix_and
   (.i_x (xdn_7),
    .i_y (r_51),
    .o_z (xar_51));



// ~xd_7 & r_52
lix_and
  #(.W (32))
  u246_lix_and
   (.i_x (xdn_7),
    .i_y (r_52),
    .o_z (xar_52));



// ~xd_7 & r_53
lix_and
  #(.W (32))
  u247_lix_and
   (.i_x (xdn_7),
    .i_y (r_53),
    .o_z (xar_53));



// ~xd_7 & r_54
lix_and
  #(.W (32))
  u248_lix_and
   (.i_x (xdn_7),
    .i_y (r_54),
    .o_z (xar_54));



// ~xd_7 & r_55
lix_and
  #(.W (32))
  u249_lix_and
   (.i_x (xdn_7),
    .i_y (r_55),
    .o_z (xar_55));



// delay ~xd_0 & r_0
lix_reg
  #(.W (32))
  u250_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_0),
    .o_z    (u_0));



// delay ~xd_1 & r_1
lix_reg
  #(.W (32))
  u251_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_1),
    .o_z    (u_1));



// delay ~xd_2 & r_2
lix_reg
  #(.W (32))
  u252_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_2),
    .o_z    (u_2));



// delay ~xd_3 & r_3
lix_reg
  #(.W (32))
  u253_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_3),
    .o_z    (u_3));



// delay ~xd_4 & r_4
lix_reg
  #(.W (32))
  u254_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_4),
    .o_z    (u_4));



// delay ~xd_5 & r_5
lix_reg
  #(.W (32))
  u255_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_5),
    .o_z    (u_5));



// delay ~xd_6 & r_6
lix_reg
  #(.W (32))
  u256_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_6),
    .o_z    (u_6));



// delay ~xd_7 & r_7
lix_reg
  #(.W (32))
  u257_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_7),
    .o_z    (u_7));



// delay ~xd_8 & r_8
lix_reg
  #(.W (32))
  u258_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_8),
    .o_z    (u_8));



// delay ~xd_9 & r_9
lix_reg
  #(.W (32))
  u259_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_9),
    .o_z    (u_9));



// delay ~xd_10 & r_10
lix_reg
  #(.W (32))
  u260_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_10),
    .o_z    (u_10));



// delay ~xd_11 & r_11
lix_reg
  #(.W (32))
  u261_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_11),
    .o_z    (u_11));



// delay ~xd_12 & r_12
lix_reg
  #(.W (32))
  u262_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_12),
    .o_z    (u_12));



// delay ~xd_13 & r_13
lix_reg
  #(.W (32))
  u263_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_13),
    .o_z    (u_13));



// delay ~xd_14 & r_14
lix_reg
  #(.W (32))
  u264_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_14),
    .o_z    (u_14));



// delay ~xd_15 & r_15
lix_reg
  #(.W (32))
  u265_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_15),
    .o_z    (u_15));



// delay ~xd_16 & r_16
lix_reg
  #(.W (32))
  u266_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_16),
    .o_z    (u_16));



// delay ~xd_17 & r_17
lix_reg
  #(.W (32))
  u267_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_17),
    .o_z    (u_17));



// delay ~xd_18 & r_18
lix_reg
  #(.W (32))
  u268_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_18),
    .o_z    (u_18));



// delay ~xd_19 & r_19
lix_reg
  #(.W (32))
  u269_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_19),
    .o_z    (u_19));



// delay ~xd_20 & r_20
lix_reg
  #(.W (32))
  u270_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_20),
    .o_z    (u_20));



// delay ~xd_21 & r_21
lix_reg
  #(.W (32))
  u271_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_21),
    .o_z    (u_21));



// delay ~xd_22 & r_22
lix_reg
  #(.W (32))
  u272_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_22),
    .o_z    (u_22));



// delay ~xd_23 & r_23
lix_reg
  #(.W (32))
  u273_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_23),
    .o_z    (u_23));



// delay ~xd_24 & r_24
lix_reg
  #(.W (32))
  u274_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_24),
    .o_z    (u_24));



// delay ~xd_25 & r_25
lix_reg
  #(.W (32))
  u275_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_25),
    .o_z    (u_25));



// delay ~xd_26 & r_26
lix_reg
  #(.W (32))
  u276_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_26),
    .o_z    (u_26));



// delay ~xd_27 & r_27
lix_reg
  #(.W (32))
  u277_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_27),
    .o_z    (u_27));



// delay ~xd_28 & r_28
lix_reg
  #(.W (32))
  u278_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_28),
    .o_z    (u_28));



// delay ~xd_29 & r_29
lix_reg
  #(.W (32))
  u279_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_29),
    .o_z    (u_29));



// delay ~xd_30 & r_30
lix_reg
  #(.W (32))
  u280_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_30),
    .o_z    (u_30));



// delay ~xd_31 & r_31
lix_reg
  #(.W (32))
  u281_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_31),
    .o_z    (u_31));



// delay ~xd_32 & r_32
lix_reg
  #(.W (32))
  u282_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_32),
    .o_z    (u_32));



// delay ~xd_33 & r_33
lix_reg
  #(.W (32))
  u283_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_33),
    .o_z    (u_33));



// delay ~xd_34 & r_34
lix_reg
  #(.W (32))
  u284_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_34),
    .o_z    (u_34));



// delay ~xd_35 & r_35
lix_reg
  #(.W (32))
  u285_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_35),
    .o_z    (u_35));



// delay ~xd_36 & r_36
lix_reg
  #(.W (32))
  u286_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_36),
    .o_z    (u_36));



// delay ~xd_37 & r_37
lix_reg
  #(.W (32))
  u287_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_37),
    .o_z    (u_37));



// delay ~xd_38 & r_38
lix_reg
  #(.W (32))
  u288_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_38),
    .o_z    (u_38));



// delay ~xd_39 & r_39
lix_reg
  #(.W (32))
  u289_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_39),
    .o_z    (u_39));



// delay ~xd_40 & r_40
lix_reg
  #(.W (32))
  u290_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_40),
    .o_z    (u_40));



// delay ~xd_41 & r_41
lix_reg
  #(.W (32))
  u291_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_41),
    .o_z    (u_41));



// delay ~xd_42 & r_42
lix_reg
  #(.W (32))
  u292_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_42),
    .o_z    (u_42));



// delay ~xd_43 & r_43
lix_reg
  #(.W (32))
  u293_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_43),
    .o_z    (u_43));



// delay ~xd_44 & r_44
lix_reg
  #(.W (32))
  u294_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_44),
    .o_z    (u_44));



// delay ~xd_45 & r_45
lix_reg
  #(.W (32))
  u295_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_45),
    .o_z    (u_45));



// delay ~xd_46 & r_46
lix_reg
  #(.W (32))
  u296_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_46),
    .o_z    (u_46));



// delay ~xd_47 & r_47
lix_reg
  #(.W (32))
  u297_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_47),
    .o_z    (u_47));



// delay ~xd_48 & r_48
lix_reg
  #(.W (32))
  u298_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_48),
    .o_z    (u_48));



// delay ~xd_49 & r_49
lix_reg
  #(.W (32))
  u299_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_49),
    .o_z    (u_49));



// delay ~xd_50 & r_50
lix_reg
  #(.W (32))
  u300_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_50),
    .o_z    (u_50));



// delay ~xd_51 & r_51
lix_reg
  #(.W (32))
  u301_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_51),
    .o_z    (u_51));



// delay ~xd_52 & r_52
lix_reg
  #(.W (32))
  u302_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_52),
    .o_z    (u_52));



// delay ~xd_53 & r_53
lix_reg
  #(.W (32))
  u303_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_53),
    .o_z    (u_53));



// delay ~xd_54 & r_54
lix_reg
  #(.W (32))
  u304_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_54),
    .o_z    (u_54));



// delay ~xd_55 & r_55
lix_reg
  #(.W (32))
  u305_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xar_55),
    .o_z    (u_55));



// xd_0 & yd_0
lix_and
  #(.W (32))
  u306_lix_and
   (.i_x (xd_0),
    .i_y (yd_0),
    .o_z (xay_0));



// xd_1 & yd_1
lix_and
  #(.W (32))
  u307_lix_and
   (.i_x (xd_1),
    .i_y (yd_1),
    .o_z (xay_1));



// xd_2 & yd_2
lix_and
  #(.W (32))
  u308_lix_and
   (.i_x (xd_2),
    .i_y (yd_2),
    .o_z (xay_2));



// xd_3 & yd_3
lix_and
  #(.W (32))
  u309_lix_and
   (.i_x (xd_3),
    .i_y (yd_3),
    .o_z (xay_3));



// xd_4 & yd_4
lix_and
  #(.W (32))
  u310_lix_and
   (.i_x (xd_4),
    .i_y (yd_4),
    .o_z (xay_4));



// xd_5 & yd_5
lix_and
  #(.W (32))
  u311_lix_and
   (.i_x (xd_5),
    .i_y (yd_5),
    .o_z (xay_5));



// xd_6 & yd_6
lix_and
  #(.W (32))
  u312_lix_and
   (.i_x (xd_6),
    .i_y (yd_6),
    .o_z (xay_6));



// xd_7 & yd_7
lix_and
  #(.W (32))
  u313_lix_and
   (.i_x (xd_7),
    .i_y (yd_7),
    .o_z (xay_7));



// delay xd_0 & yd_0
lix_reg
  #(.W (32))
  u314_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_0),
    .o_z    (k_0));



// delay xd_1 & yd_1
lix_reg
  #(.W (32))
  u315_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_1),
    .o_z    (k_1));



// delay xd_2 & yd_2
lix_reg
  #(.W (32))
  u316_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_2),
    .o_z    (k_2));



// delay xd_3 & yd_3
lix_reg
  #(.W (32))
  u317_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_3),
    .o_z    (k_3));



// delay xd_4 & yd_4
lix_reg
  #(.W (32))
  u318_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_4),
    .o_z    (k_4));



// delay xd_5 & yd_5
lix_reg
  #(.W (32))
  u319_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_5),
    .o_z    (k_5));



// delay xd_6 & yd_6
lix_reg
  #(.W (32))
  u320_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_6),
    .o_z    (k_6));



// delay xd_7 & yd_7
lix_reg
  #(.W (32))
  u321_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xay_7),
    .o_z    (k_7));



// xd_0 & v_0
lix_and
  #(.W (32))
  u322_lix_and
   (.i_x (xd_0),
    .i_y (v_0),
    .o_z (xav_0));



// xd_0 & v_1
lix_and
  #(.W (32))
  u323_lix_and
   (.i_x (xd_0),
    .i_y (v_1),
    .o_z (xav_1));



// xd_0 & v_2
lix_and
  #(.W (32))
  u324_lix_and
   (.i_x (xd_0),
    .i_y (v_2),
    .o_z (xav_2));



// xd_0 & v_3
lix_and
  #(.W (32))
  u325_lix_and
   (.i_x (xd_0),
    .i_y (v_3),
    .o_z (xav_3));



// xd_0 & v_4
lix_and
  #(.W (32))
  u326_lix_and
   (.i_x (xd_0),
    .i_y (v_4),
    .o_z (xav_4));



// xd_0 & v_5
lix_and
  #(.W (32))
  u327_lix_and
   (.i_x (xd_0),
    .i_y (v_5),
    .o_z (xav_5));



// xd_0 & v_6
lix_and
  #(.W (32))
  u328_lix_and
   (.i_x (xd_0),
    .i_y (v_6),
    .o_z (xav_6));



// xd_1 & v_7
lix_and
  #(.W (32))
  u329_lix_and
   (.i_x (xd_1),
    .i_y (v_7),
    .o_z (xav_7));



// xd_1 & v_8
lix_and
  #(.W (32))
  u330_lix_and
   (.i_x (xd_1),
    .i_y (v_8),
    .o_z (xav_8));



// xd_1 & v_9
lix_and
  #(.W (32))
  u331_lix_and
   (.i_x (xd_1),
    .i_y (v_9),
    .o_z (xav_9));



// xd_1 & v_10
lix_and
  #(.W (32))
  u332_lix_and
   (.i_x (xd_1),
    .i_y (v_10),
    .o_z (xav_10));



// xd_1 & v_11
lix_and
  #(.W (32))
  u333_lix_and
   (.i_x (xd_1),
    .i_y (v_11),
    .o_z (xav_11));



// xd_1 & v_12
lix_and
  #(.W (32))
  u334_lix_and
   (.i_x (xd_1),
    .i_y (v_12),
    .o_z (xav_12));



// xd_1 & v_13
lix_and
  #(.W (32))
  u335_lix_and
   (.i_x (xd_1),
    .i_y (v_13),
    .o_z (xav_13));



// xd_2 & v_14
lix_and
  #(.W (32))
  u336_lix_and
   (.i_x (xd_2),
    .i_y (v_14),
    .o_z (xav_14));



// xd_2 & v_15
lix_and
  #(.W (32))
  u337_lix_and
   (.i_x (xd_2),
    .i_y (v_15),
    .o_z (xav_15));



// xd_2 & v_16
lix_and
  #(.W (32))
  u338_lix_and
   (.i_x (xd_2),
    .i_y (v_16),
    .o_z (xav_16));



// xd_2 & v_17
lix_and
  #(.W (32))
  u339_lix_and
   (.i_x (xd_2),
    .i_y (v_17),
    .o_z (xav_17));



// xd_2 & v_18
lix_and
  #(.W (32))
  u340_lix_and
   (.i_x (xd_2),
    .i_y (v_18),
    .o_z (xav_18));



// xd_2 & v_19
lix_and
  #(.W (32))
  u341_lix_and
   (.i_x (xd_2),
    .i_y (v_19),
    .o_z (xav_19));



// xd_2 & v_20
lix_and
  #(.W (32))
  u342_lix_and
   (.i_x (xd_2),
    .i_y (v_20),
    .o_z (xav_20));



// xd_3 & v_21
lix_and
  #(.W (32))
  u343_lix_and
   (.i_x (xd_3),
    .i_y (v_21),
    .o_z (xav_21));



// xd_3 & v_22
lix_and
  #(.W (32))
  u344_lix_and
   (.i_x (xd_3),
    .i_y (v_22),
    .o_z (xav_22));



// xd_3 & v_23
lix_and
  #(.W (32))
  u345_lix_and
   (.i_x (xd_3),
    .i_y (v_23),
    .o_z (xav_23));



// xd_3 & v_24
lix_and
  #(.W (32))
  u346_lix_and
   (.i_x (xd_3),
    .i_y (v_24),
    .o_z (xav_24));



// xd_3 & v_25
lix_and
  #(.W (32))
  u347_lix_and
   (.i_x (xd_3),
    .i_y (v_25),
    .o_z (xav_25));



// xd_3 & v_26
lix_and
  #(.W (32))
  u348_lix_and
   (.i_x (xd_3),
    .i_y (v_26),
    .o_z (xav_26));



// xd_3 & v_27
lix_and
  #(.W (32))
  u349_lix_and
   (.i_x (xd_3),
    .i_y (v_27),
    .o_z (xav_27));



// xd_4 & v_28
lix_and
  #(.W (32))
  u350_lix_and
   (.i_x (xd_4),
    .i_y (v_28),
    .o_z (xav_28));



// xd_4 & v_29
lix_and
  #(.W (32))
  u351_lix_and
   (.i_x (xd_4),
    .i_y (v_29),
    .o_z (xav_29));



// xd_4 & v_30
lix_and
  #(.W (32))
  u352_lix_and
   (.i_x (xd_4),
    .i_y (v_30),
    .o_z (xav_30));



// xd_4 & v_31
lix_and
  #(.W (32))
  u353_lix_and
   (.i_x (xd_4),
    .i_y (v_31),
    .o_z (xav_31));



// xd_4 & v_32
lix_and
  #(.W (32))
  u354_lix_and
   (.i_x (xd_4),
    .i_y (v_32),
    .o_z (xav_32));



// xd_4 & v_33
lix_and
  #(.W (32))
  u355_lix_and
   (.i_x (xd_4),
    .i_y (v_33),
    .o_z (xav_33));



// xd_4 & v_34
lix_and
  #(.W (32))
  u356_lix_and
   (.i_x (xd_4),
    .i_y (v_34),
    .o_z (xav_34));



// xd_5 & v_35
lix_and
  #(.W (32))
  u357_lix_and
   (.i_x (xd_5),
    .i_y (v_35),
    .o_z (xav_35));



// xd_5 & v_36
lix_and
  #(.W (32))
  u358_lix_and
   (.i_x (xd_5),
    .i_y (v_36),
    .o_z (xav_36));



// xd_5 & v_37
lix_and
  #(.W (32))
  u359_lix_and
   (.i_x (xd_5),
    .i_y (v_37),
    .o_z (xav_37));



// xd_5 & v_38
lix_and
  #(.W (32))
  u360_lix_and
   (.i_x (xd_5),
    .i_y (v_38),
    .o_z (xav_38));



// xd_5 & v_39
lix_and
  #(.W (32))
  u361_lix_and
   (.i_x (xd_5),
    .i_y (v_39),
    .o_z (xav_39));



// xd_5 & v_40
lix_and
  #(.W (32))
  u362_lix_and
   (.i_x (xd_5),
    .i_y (v_40),
    .o_z (xav_40));



// xd_5 & v_41
lix_and
  #(.W (32))
  u363_lix_and
   (.i_x (xd_5),
    .i_y (v_41),
    .o_z (xav_41));



// xd_6 & v_42
lix_and
  #(.W (32))
  u364_lix_and
   (.i_x (xd_6),
    .i_y (v_42),
    .o_z (xav_42));



// xd_6 & v_43
lix_and
  #(.W (32))
  u365_lix_and
   (.i_x (xd_6),
    .i_y (v_43),
    .o_z (xav_43));



// xd_6 & v_44
lix_and
  #(.W (32))
  u366_lix_and
   (.i_x (xd_6),
    .i_y (v_44),
    .o_z (xav_44));



// xd_6 & v_45
lix_and
  #(.W (32))
  u367_lix_and
   (.i_x (xd_6),
    .i_y (v_45),
    .o_z (xav_45));



// xd_6 & v_46
lix_and
  #(.W (32))
  u368_lix_and
   (.i_x (xd_6),
    .i_y (v_46),
    .o_z (xav_46));



// xd_6 & v_47
lix_and
  #(.W (32))
  u369_lix_and
   (.i_x (xd_6),
    .i_y (v_47),
    .o_z (xav_47));



// xd_6 & v_48
lix_and
  #(.W (32))
  u370_lix_and
   (.i_x (xd_6),
    .i_y (v_48),
    .o_z (xav_48));



// xd_7 & v_49
lix_and
  #(.W (32))
  u371_lix_and
   (.i_x (xd_7),
    .i_y (v_49),
    .o_z (xav_49));



// xd_7 & v_50
lix_and
  #(.W (32))
  u372_lix_and
   (.i_x (xd_7),
    .i_y (v_50),
    .o_z (xav_50));



// xd_7 & v_51
lix_and
  #(.W (32))
  u373_lix_and
   (.i_x (xd_7),
    .i_y (v_51),
    .o_z (xav_51));



// xd_7 & v_52
lix_and
  #(.W (32))
  u374_lix_and
   (.i_x (xd_7),
    .i_y (v_52),
    .o_z (xav_52));



// xd_7 & v_53
lix_and
  #(.W (32))
  u375_lix_and
   (.i_x (xd_7),
    .i_y (v_53),
    .o_z (xav_53));



// xd_7 & v_54
lix_and
  #(.W (32))
  u376_lix_and
   (.i_x (xd_7),
    .i_y (v_54),
    .o_z (xav_54));



// xd_7 & v_55
lix_and
  #(.W (32))
  u377_lix_and
   (.i_x (xd_7),
    .i_y (v_55),
    .o_z (xav_55));



// delay xd_0 & v_0
lix_reg
  #(.W (32))
  u378_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_0),
    .o_z    (t_0));



// delay xd_1 & v_1
lix_reg
  #(.W (32))
  u379_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_1),
    .o_z    (t_1));



// delay xd_2 & v_2
lix_reg
  #(.W (32))
  u380_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_2),
    .o_z    (t_2));



// delay xd_3 & v_3
lix_reg
  #(.W (32))
  u381_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_3),
    .o_z    (t_3));



// delay xd_4 & v_4
lix_reg
  #(.W (32))
  u382_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_4),
    .o_z    (t_4));



// delay xd_5 & v_5
lix_reg
  #(.W (32))
  u383_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_5),
    .o_z    (t_5));



// delay xd_6 & v_6
lix_reg
  #(.W (32))
  u384_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_6),
    .o_z    (t_6));



// delay xd_7 & v_7
lix_reg
  #(.W (32))
  u385_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_7),
    .o_z    (t_7));



// delay xd_8 & v_8
lix_reg
  #(.W (32))
  u386_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_8),
    .o_z    (t_8));



// delay xd_9 & v_9
lix_reg
  #(.W (32))
  u387_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_9),
    .o_z    (t_9));



// delay xd_10 & v_10
lix_reg
  #(.W (32))
  u388_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_10),
    .o_z    (t_10));



// delay xd_11 & v_11
lix_reg
  #(.W (32))
  u389_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_11),
    .o_z    (t_11));



// delay xd_12 & v_12
lix_reg
  #(.W (32))
  u390_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_12),
    .o_z    (t_12));



// delay xd_13 & v_13
lix_reg
  #(.W (32))
  u391_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_13),
    .o_z    (t_13));



// delay xd_14 & v_14
lix_reg
  #(.W (32))
  u392_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_14),
    .o_z    (t_14));



// delay xd_15 & v_15
lix_reg
  #(.W (32))
  u393_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_15),
    .o_z    (t_15));



// delay xd_16 & v_16
lix_reg
  #(.W (32))
  u394_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_16),
    .o_z    (t_16));



// delay xd_17 & v_17
lix_reg
  #(.W (32))
  u395_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_17),
    .o_z    (t_17));



// delay xd_18 & v_18
lix_reg
  #(.W (32))
  u396_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_18),
    .o_z    (t_18));



// delay xd_19 & v_19
lix_reg
  #(.W (32))
  u397_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_19),
    .o_z    (t_19));



// delay xd_20 & v_20
lix_reg
  #(.W (32))
  u398_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_20),
    .o_z    (t_20));



// delay xd_21 & v_21
lix_reg
  #(.W (32))
  u399_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_21),
    .o_z    (t_21));



// delay xd_22 & v_22
lix_reg
  #(.W (32))
  u400_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_22),
    .o_z    (t_22));



// delay xd_23 & v_23
lix_reg
  #(.W (32))
  u401_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_23),
    .o_z    (t_23));



// delay xd_24 & v_24
lix_reg
  #(.W (32))
  u402_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_24),
    .o_z    (t_24));



// delay xd_25 & v_25
lix_reg
  #(.W (32))
  u403_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_25),
    .o_z    (t_25));



// delay xd_26 & v_26
lix_reg
  #(.W (32))
  u404_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_26),
    .o_z    (t_26));



// delay xd_27 & v_27
lix_reg
  #(.W (32))
  u405_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_27),
    .o_z    (t_27));



// delay xd_28 & v_28
lix_reg
  #(.W (32))
  u406_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_28),
    .o_z    (t_28));



// delay xd_29 & v_29
lix_reg
  #(.W (32))
  u407_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_29),
    .o_z    (t_29));



// delay xd_30 & v_30
lix_reg
  #(.W (32))
  u408_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_30),
    .o_z    (t_30));



// delay xd_31 & v_31
lix_reg
  #(.W (32))
  u409_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_31),
    .o_z    (t_31));



// delay xd_32 & v_32
lix_reg
  #(.W (32))
  u410_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_32),
    .o_z    (t_32));



// delay xd_33 & v_33
lix_reg
  #(.W (32))
  u411_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_33),
    .o_z    (t_33));



// delay xd_34 & v_34
lix_reg
  #(.W (32))
  u412_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_34),
    .o_z    (t_34));



// delay xd_35 & v_35
lix_reg
  #(.W (32))
  u413_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_35),
    .o_z    (t_35));



// delay xd_36 & v_36
lix_reg
  #(.W (32))
  u414_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_36),
    .o_z    (t_36));



// delay xd_37 & v_37
lix_reg
  #(.W (32))
  u415_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_37),
    .o_z    (t_37));



// delay xd_38 & v_38
lix_reg
  #(.W (32))
  u416_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_38),
    .o_z    (t_38));



// delay xd_39 & v_39
lix_reg
  #(.W (32))
  u417_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_39),
    .o_z    (t_39));



// delay xd_40 & v_40
lix_reg
  #(.W (32))
  u418_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_40),
    .o_z    (t_40));



// delay xd_41 & v_41
lix_reg
  #(.W (32))
  u419_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_41),
    .o_z    (t_41));



// delay xd_42 & v_42
lix_reg
  #(.W (32))
  u420_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_42),
    .o_z    (t_42));



// delay xd_43 & v_43
lix_reg
  #(.W (32))
  u421_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_43),
    .o_z    (t_43));



// delay xd_44 & v_44
lix_reg
  #(.W (32))
  u422_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_44),
    .o_z    (t_44));



// delay xd_45 & v_45
lix_reg
  #(.W (32))
  u423_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_45),
    .o_z    (t_45));



// delay xd_46 & v_46
lix_reg
  #(.W (32))
  u424_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_46),
    .o_z    (t_46));



// delay xd_47 & v_47
lix_reg
  #(.W (32))
  u425_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_47),
    .o_z    (t_47));



// delay xd_48 & v_48
lix_reg
  #(.W (32))
  u426_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_48),
    .o_z    (t_48));



// delay xd_49 & v_49
lix_reg
  #(.W (32))
  u427_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_49),
    .o_z    (t_49));



// delay xd_50 & v_50
lix_reg
  #(.W (32))
  u428_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_50),
    .o_z    (t_50));



// delay xd_51 & v_51
lix_reg
  #(.W (32))
  u429_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_51),
    .o_z    (t_51));



// delay xd_52 & v_52
lix_reg
  #(.W (32))
  u430_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_52),
    .o_z    (t_52));



// delay xd_53 & v_53
lix_reg
  #(.W (32))
  u431_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_53),
    .o_z    (t_53));



// delay xd_54 & v_54
lix_reg
  #(.W (32))
  u432_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_54),
    .o_z    (t_54));



// delay xd_55 & v_55
lix_reg
  #(.W (32))
  u433_lix_reg
   (.clk_i  (clk_i),
    .rst_ni (rst_ni),
    .i_vld  (vldd1),
    .i_en   (i_rvld),
    .i_x    (xav_55),
    .o_z    (t_55));



// u_0 ^ t_0
lix_xor
  #(.W (32))
  u434_lix_xor
   (.i_x (u_0),
    .i_y (t_0),
    .o_z (z_0));



// u_1 ^ t_1
lix_xor
  #(.W (32))
  u435_lix_xor
   (.i_x (u_1),
    .i_y (t_1),
    .o_z (z_1));



// u_2 ^ t_2
lix_xor
  #(.W (32))
  u436_lix_xor
   (.i_x (u_2),
    .i_y (t_2),
    .o_z (z_2));



// u_3 ^ t_3
lix_xor
  #(.W (32))
  u437_lix_xor
   (.i_x (u_3),
    .i_y (t_3),
    .o_z (z_3));



// u_4 ^ t_4
lix_xor
  #(.W (32))
  u438_lix_xor
   (.i_x (u_4),
    .i_y (t_4),
    .o_z (z_4));



// u_5 ^ t_5
lix_xor
  #(.W (32))
  u439_lix_xor
   (.i_x (u_5),
    .i_y (t_5),
    .o_z (z_5));



// u_6 ^ t_6
lix_xor
  #(.W (32))
  u440_lix_xor
   (.i_x (u_6),
    .i_y (t_6),
    .o_z (z_6));



// u_7 ^ t_7
lix_xor
  #(.W (32))
  u441_lix_xor
   (.i_x (u_7),
    .i_y (t_7),
    .o_z (z_7));



// u_8 ^ t_8
lix_xor
  #(.W (32))
  u442_lix_xor
   (.i_x (u_8),
    .i_y (t_8),
    .o_z (z_8));



// u_9 ^ t_9
lix_xor
  #(.W (32))
  u443_lix_xor
   (.i_x (u_9),
    .i_y (t_9),
    .o_z (z_9));



// u_10 ^ t_10
lix_xor
  #(.W (32))
  u444_lix_xor
   (.i_x (u_10),
    .i_y (t_10),
    .o_z (z_10));



// u_11 ^ t_11
lix_xor
  #(.W (32))
  u445_lix_xor
   (.i_x (u_11),
    .i_y (t_11),
    .o_z (z_11));



// u_12 ^ t_12
lix_xor
  #(.W (32))
  u446_lix_xor
   (.i_x (u_12),
    .i_y (t_12),
    .o_z (z_12));



// u_13 ^ t_13
lix_xor
  #(.W (32))
  u447_lix_xor
   (.i_x (u_13),
    .i_y (t_13),
    .o_z (z_13));



// u_14 ^ t_14
lix_xor
  #(.W (32))
  u448_lix_xor
   (.i_x (u_14),
    .i_y (t_14),
    .o_z (z_14));



// u_15 ^ t_15
lix_xor
  #(.W (32))
  u449_lix_xor
   (.i_x (u_15),
    .i_y (t_15),
    .o_z (z_15));



// u_16 ^ t_16
lix_xor
  #(.W (32))
  u450_lix_xor
   (.i_x (u_16),
    .i_y (t_16),
    .o_z (z_16));



// u_17 ^ t_17
lix_xor
  #(.W (32))
  u451_lix_xor
   (.i_x (u_17),
    .i_y (t_17),
    .o_z (z_17));



// u_18 ^ t_18
lix_xor
  #(.W (32))
  u452_lix_xor
   (.i_x (u_18),
    .i_y (t_18),
    .o_z (z_18));



// u_19 ^ t_19
lix_xor
  #(.W (32))
  u453_lix_xor
   (.i_x (u_19),
    .i_y (t_19),
    .o_z (z_19));



// u_20 ^ t_20
lix_xor
  #(.W (32))
  u454_lix_xor
   (.i_x (u_20),
    .i_y (t_20),
    .o_z (z_20));



// u_21 ^ t_21
lix_xor
  #(.W (32))
  u455_lix_xor
   (.i_x (u_21),
    .i_y (t_21),
    .o_z (z_21));



// u_22 ^ t_22
lix_xor
  #(.W (32))
  u456_lix_xor
   (.i_x (u_22),
    .i_y (t_22),
    .o_z (z_22));



// u_23 ^ t_23
lix_xor
  #(.W (32))
  u457_lix_xor
   (.i_x (u_23),
    .i_y (t_23),
    .o_z (z_23));



// u_24 ^ t_24
lix_xor
  #(.W (32))
  u458_lix_xor
   (.i_x (u_24),
    .i_y (t_24),
    .o_z (z_24));



// u_25 ^ t_25
lix_xor
  #(.W (32))
  u459_lix_xor
   (.i_x (u_25),
    .i_y (t_25),
    .o_z (z_25));



// u_26 ^ t_26
lix_xor
  #(.W (32))
  u460_lix_xor
   (.i_x (u_26),
    .i_y (t_26),
    .o_z (z_26));



// u_27 ^ t_27
lix_xor
  #(.W (32))
  u461_lix_xor
   (.i_x (u_27),
    .i_y (t_27),
    .o_z (z_27));



// u_28 ^ t_28
lix_xor
  #(.W (32))
  u462_lix_xor
   (.i_x (u_28),
    .i_y (t_28),
    .o_z (z_28));



// u_29 ^ t_29
lix_xor
  #(.W (32))
  u463_lix_xor
   (.i_x (u_29),
    .i_y (t_29),
    .o_z (z_29));



// u_30 ^ t_30
lix_xor
  #(.W (32))
  u464_lix_xor
   (.i_x (u_30),
    .i_y (t_30),
    .o_z (z_30));



// u_31 ^ t_31
lix_xor
  #(.W (32))
  u465_lix_xor
   (.i_x (u_31),
    .i_y (t_31),
    .o_z (z_31));



// u_32 ^ t_32
lix_xor
  #(.W (32))
  u466_lix_xor
   (.i_x (u_32),
    .i_y (t_32),
    .o_z (z_32));



// u_33 ^ t_33
lix_xor
  #(.W (32))
  u467_lix_xor
   (.i_x (u_33),
    .i_y (t_33),
    .o_z (z_33));



// u_34 ^ t_34
lix_xor
  #(.W (32))
  u468_lix_xor
   (.i_x (u_34),
    .i_y (t_34),
    .o_z (z_34));



// u_35 ^ t_35
lix_xor
  #(.W (32))
  u469_lix_xor
   (.i_x (u_35),
    .i_y (t_35),
    .o_z (z_35));



// u_36 ^ t_36
lix_xor
  #(.W (32))
  u470_lix_xor
   (.i_x (u_36),
    .i_y (t_36),
    .o_z (z_36));



// u_37 ^ t_37
lix_xor
  #(.W (32))
  u471_lix_xor
   (.i_x (u_37),
    .i_y (t_37),
    .o_z (z_37));



// u_38 ^ t_38
lix_xor
  #(.W (32))
  u472_lix_xor
   (.i_x (u_38),
    .i_y (t_38),
    .o_z (z_38));



// u_39 ^ t_39
lix_xor
  #(.W (32))
  u473_lix_xor
   (.i_x (u_39),
    .i_y (t_39),
    .o_z (z_39));



// u_40 ^ t_40
lix_xor
  #(.W (32))
  u474_lix_xor
   (.i_x (u_40),
    .i_y (t_40),
    .o_z (z_40));



// u_41 ^ t_41
lix_xor
  #(.W (32))
  u475_lix_xor
   (.i_x (u_41),
    .i_y (t_41),
    .o_z (z_41));



// u_42 ^ t_42
lix_xor
  #(.W (32))
  u476_lix_xor
   (.i_x (u_42),
    .i_y (t_42),
    .o_z (z_42));



// u_43 ^ t_43
lix_xor
  #(.W (32))
  u477_lix_xor
   (.i_x (u_43),
    .i_y (t_43),
    .o_z (z_43));



// u_44 ^ t_44
lix_xor
  #(.W (32))
  u478_lix_xor
   (.i_x (u_44),
    .i_y (t_44),
    .o_z (z_44));



// u_45 ^ t_45
lix_xor
  #(.W (32))
  u479_lix_xor
   (.i_x (u_45),
    .i_y (t_45),
    .o_z (z_45));



// u_46 ^ t_46
lix_xor
  #(.W (32))
  u480_lix_xor
   (.i_x (u_46),
    .i_y (t_46),
    .o_z (z_46));



// u_47 ^ t_47
lix_xor
  #(.W (32))
  u481_lix_xor
   (.i_x (u_47),
    .i_y (t_47),
    .o_z (z_47));



// u_48 ^ t_48
lix_xor
  #(.W (32))
  u482_lix_xor
   (.i_x (u_48),
    .i_y (t_48),
    .o_z (z_48));



// u_49 ^ t_49
lix_xor
  #(.W (32))
  u483_lix_xor
   (.i_x (u_49),
    .i_y (t_49),
    .o_z (z_49));



// u_50 ^ t_50
lix_xor
  #(.W (32))
  u484_lix_xor
   (.i_x (u_50),
    .i_y (t_50),
    .o_z (z_50));



// u_51 ^ t_51
lix_xor
  #(.W (32))
  u485_lix_xor
   (.i_x (u_51),
    .i_y (t_51),
    .o_z (z_51));



// u_52 ^ t_52
lix_xor
  #(.W (32))
  u486_lix_xor
   (.i_x (u_52),
    .i_y (t_52),
    .o_z (z_52));



// u_53 ^ t_53
lix_xor
  #(.W (32))
  u487_lix_xor
   (.i_x (u_53),
    .i_y (t_53),
    .o_z (z_53));



// u_54 ^ t_54
lix_xor
  #(.W (32))
  u488_lix_xor
   (.i_x (u_54),
    .i_y (t_54),
    .o_z (z_54));



// u_55 ^ t_55
lix_xor
  #(.W (32))
  u489_lix_xor
   (.i_x (u_55),
    .i_y (t_55),
    .o_z (z_55));



// z_1 ^ z_0
lix_xor
  #(.W (32))
  u490_lix_xor
   (.i_x (z_0),
    .i_y (z_1),
    .o_z (zxz_0));



// z_2 ^ zxz_0
lix_xor
  #(.W (32))
  u491_lix_xor
   (.i_x (z_2),
    .i_y (zxz_0),
    .o_z (zxz_1));



// z_3 ^ zxz_1
lix_xor
  #(.W (32))
  u492_lix_xor
   (.i_x (z_3),
    .i_y (zxz_1),
    .o_z (zxz_2));



// z_4 ^ zxz_2
lix_xor
  #(.W (32))
  u493_lix_xor
   (.i_x (z_4),
    .i_y (zxz_2),
    .o_z (zxz_3));



// z_5 ^ zxz_3
lix_xor
  #(.W (32))
  u494_lix_xor
   (.i_x (z_5),
    .i_y (zxz_3),
    .o_z (zxz_4));



// z_6 ^ zxz_4
lix_xor
  #(.W (32))
  u495_lix_xor
   (.i_x (z_6),
    .i_y (zxz_4),
    .o_z (zxz_5));



// z_8 ^ z_7
lix_xor
  #(.W (32))
  u496_lix_xor
   (.i_x (z_7),
    .i_y (z_8),
    .o_z (zxz_6));



// z_9 ^ zxz_6
lix_xor
  #(.W (32))
  u497_lix_xor
   (.i_x (z_9),
    .i_y (zxz_6),
    .o_z (zxz_7));



// z_10 ^ zxz_7
lix_xor
  #(.W (32))
  u498_lix_xor
   (.i_x (z_10),
    .i_y (zxz_7),
    .o_z (zxz_8));



// z_11 ^ zxz_8
lix_xor
  #(.W (32))
  u499_lix_xor
   (.i_x (z_11),
    .i_y (zxz_8),
    .o_z (zxz_9));



// z_12 ^ zxz_9
lix_xor
  #(.W (32))
  u500_lix_xor
   (.i_x (z_12),
    .i_y (zxz_9),
    .o_z (zxz_10));



// z_13 ^ zxz_10
lix_xor
  #(.W (32))
  u501_lix_xor
   (.i_x (z_13),
    .i_y (zxz_10),
    .o_z (zxz_11));



// z_15 ^ z_14
lix_xor
  #(.W (32))
  u502_lix_xor
   (.i_x (z_14),
    .i_y (z_15),
    .o_z (zxz_12));



// z_16 ^ zxz_12
lix_xor
  #(.W (32))
  u503_lix_xor
   (.i_x (z_16),
    .i_y (zxz_12),
    .o_z (zxz_13));



// z_17 ^ zxz_13
lix_xor
  #(.W (32))
  u504_lix_xor
   (.i_x (z_17),
    .i_y (zxz_13),
    .o_z (zxz_14));



// z_18 ^ zxz_14
lix_xor
  #(.W (32))
  u505_lix_xor
   (.i_x (z_18),
    .i_y (zxz_14),
    .o_z (zxz_15));



// z_19 ^ zxz_15
lix_xor
  #(.W (32))
  u506_lix_xor
   (.i_x (z_19),
    .i_y (zxz_15),
    .o_z (zxz_16));



// z_20 ^ zxz_16
lix_xor
  #(.W (32))
  u507_lix_xor
   (.i_x (z_20),
    .i_y (zxz_16),
    .o_z (zxz_17));



// z_22 ^ z_21
lix_xor
  #(.W (32))
  u508_lix_xor
   (.i_x (z_21),
    .i_y (z_22),
    .o_z (zxz_18));



// z_23 ^ zxz_18
lix_xor
  #(.W (32))
  u509_lix_xor
   (.i_x (z_23),
    .i_y (zxz_18),
    .o_z (zxz_19));



// z_24 ^ zxz_19
lix_xor
  #(.W (32))
  u510_lix_xor
   (.i_x (z_24),
    .i_y (zxz_19),
    .o_z (zxz_20));



// z_25 ^ zxz_20
lix_xor
  #(.W (32))
  u511_lix_xor
   (.i_x (z_25),
    .i_y (zxz_20),
    .o_z (zxz_21));



// z_26 ^ zxz_21
lix_xor
  #(.W (32))
  u512_lix_xor
   (.i_x (z_26),
    .i_y (zxz_21),
    .o_z (zxz_22));



// z_27 ^ zxz_22
lix_xor
  #(.W (32))
  u513_lix_xor
   (.i_x (z_27),
    .i_y (zxz_22),
    .o_z (zxz_23));



// z_29 ^ z_28
lix_xor
  #(.W (32))
  u514_lix_xor
   (.i_x (z_28),
    .i_y (z_29),
    .o_z (zxz_24));



// z_30 ^ zxz_24
lix_xor
  #(.W (32))
  u515_lix_xor
   (.i_x (z_30),
    .i_y (zxz_24),
    .o_z (zxz_25));



// z_31 ^ zxz_25
lix_xor
  #(.W (32))
  u516_lix_xor
   (.i_x (z_31),
    .i_y (zxz_25),
    .o_z (zxz_26));



// z_32 ^ zxz_26
lix_xor
  #(.W (32))
  u517_lix_xor
   (.i_x (z_32),
    .i_y (zxz_26),
    .o_z (zxz_27));



// z_33 ^ zxz_27
lix_xor
  #(.W (32))
  u518_lix_xor
   (.i_x (z_33),
    .i_y (zxz_27),
    .o_z (zxz_28));



// z_34 ^ zxz_28
lix_xor
  #(.W (32))
  u519_lix_xor
   (.i_x (z_34),
    .i_y (zxz_28),
    .o_z (zxz_29));



// z_36 ^ z_35
lix_xor
  #(.W (32))
  u520_lix_xor
   (.i_x (z_35),
    .i_y (z_36),
    .o_z (zxz_30));



// z_37 ^ zxz_30
lix_xor
  #(.W (32))
  u521_lix_xor
   (.i_x (z_37),
    .i_y (zxz_30),
    .o_z (zxz_31));



// z_38 ^ zxz_31
lix_xor
  #(.W (32))
  u522_lix_xor
   (.i_x (z_38),
    .i_y (zxz_31),
    .o_z (zxz_32));



// z_39 ^ zxz_32
lix_xor
  #(.W (32))
  u523_lix_xor
   (.i_x (z_39),
    .i_y (zxz_32),
    .o_z (zxz_33));



// z_40 ^ zxz_33
lix_xor
  #(.W (32))
  u524_lix_xor
   (.i_x (z_40),
    .i_y (zxz_33),
    .o_z (zxz_34));



// z_41 ^ zxz_34
lix_xor
  #(.W (32))
  u525_lix_xor
   (.i_x (z_41),
    .i_y (zxz_34),
    .o_z (zxz_35));



// z_43 ^ z_42
lix_xor
  #(.W (32))
  u526_lix_xor
   (.i_x (z_42),
    .i_y (z_43),
    .o_z (zxz_36));



// z_44 ^ zxz_36
lix_xor
  #(.W (32))
  u527_lix_xor
   (.i_x (z_44),
    .i_y (zxz_36),
    .o_z (zxz_37));



// z_45 ^ zxz_37
lix_xor
  #(.W (32))
  u528_lix_xor
   (.i_x (z_45),
    .i_y (zxz_37),
    .o_z (zxz_38));



// z_46 ^ zxz_38
lix_xor
  #(.W (32))
  u529_lix_xor
   (.i_x (z_46),
    .i_y (zxz_38),
    .o_z (zxz_39));



// z_47 ^ zxz_39
lix_xor
  #(.W (32))
  u530_lix_xor
   (.i_x (z_47),
    .i_y (zxz_39),
    .o_z (zxz_40));



// z_48 ^ zxz_40
lix_xor
  #(.W (32))
  u531_lix_xor
   (.i_x (z_48),
    .i_y (zxz_40),
    .o_z (zxz_41));



// z_50 ^ z_49
lix_xor
  #(.W (32))
  u532_lix_xor
   (.i_x (z_49),
    .i_y (z_50),
    .o_z (zxz_42));



// z_51 ^ zxz_42
lix_xor
  #(.W (32))
  u533_lix_xor
   (.i_x (z_51),
    .i_y (zxz_42),
    .o_z (zxz_43));



// z_52 ^ zxz_43
lix_xor
  #(.W (32))
  u534_lix_xor
   (.i_x (z_52),
    .i_y (zxz_43),
    .o_z (zxz_44));



// z_53 ^ zxz_44
lix_xor
  #(.W (32))
  u535_lix_xor
   (.i_x (z_53),
    .i_y (zxz_44),
    .o_z (zxz_45));



// z_54 ^ zxz_45
lix_xor
  #(.W (32))
  u536_lix_xor
   (.i_x (z_54),
    .i_y (zxz_45),
    .o_z (zxz_46));



// z_55 ^ zxz_46
lix_xor
  #(.W (32))
  u537_lix_xor
   (.i_x (z_55),
    .i_y (zxz_46),
    .o_z (zxz_47));



// k_0 ^ zxz_5
lix_xor
  #(.W (32))
  u538_lix_xor
   (.i_x (k_0),
    .i_y (zxz_5),
    .o_z (o_c[0+:32]));



// k_1 ^ zxz_11
lix_xor
  #(.W (32))
  u539_lix_xor
   (.i_x (k_1),
    .i_y (zxz_11),
    .o_z (o_c[32+:32]));



// k_2 ^ zxz_17
lix_xor
  #(.W (32))
  u540_lix_xor
   (.i_x (k_2),
    .i_y (zxz_17),
    .o_z (o_c[64+:32]));



// k_3 ^ zxz_23
lix_xor
  #(.W (32))
  u541_lix_xor
   (.i_x (k_3),
    .i_y (zxz_23),
    .o_z (o_c[96+:32]));



// k_4 ^ zxz_29
lix_xor
  #(.W (32))
  u542_lix_xor
   (.i_x (k_4),
    .i_y (zxz_29),
    .o_z (o_c[128+:32]));



// k_5 ^ zxz_35
lix_xor
  #(.W (32))
  u543_lix_xor
   (.i_x (k_5),
    .i_y (zxz_35),
    .o_z (o_c[160+:32]));



// k_6 ^ zxz_41
lix_xor
  #(.W (32))
  u544_lix_xor
   (.i_x (k_6),
    .i_y (zxz_41),
    .o_z (o_c[192+:32]));



// k_7 ^ zxz_47
lix_xor
  #(.W (32))
  u545_lix_xor
   (.i_x (k_7),
    .i_y (zxz_47),
    .o_z (o_c[224+:32]));



assign o_dvld = vldd2;

endmodule
